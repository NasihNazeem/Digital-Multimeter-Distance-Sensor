
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0);
		err_flag			:  OUT	STD_LOGIC
		);
END voltage2distance;

ARCHITECTURE behavior OF voltage2distance IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	1404400	)	,
(	702153	)	,
(	468071	)	,
(	351029	)	,
(	280805	)	,
(	233988	)	,
(	200548	)	,
(	175468	)	,
(	155961	)	,
(	140355	)	,
(	127587	)	,
(	116947	)	,
(	107944	)	,
(	100227	)	,
(	93539	)	,
(	87687	)	,
(	82523	)	,
(	77933	)	,
(	73827	)	,
(	70130	)	,
(	66786	)	,
(	63746	)	,
(	60971	)	,
(	58426	)	,
(	56086	)	,
(	53925	)	,
(	51924	)	,
(	50066	)	,
(	48337	)	,
(	46722	)	,
(	45212	)	,
(	43796	)	,
(	42466	)	,
(	41214	)	,
(	40034	)	,
(	38919	)	,
(	37865	)	,
(	36866	)	,
(	35918	)	,
(	35018	)	,
(	34162	)	,
(	33346	)	,
(	32568	)	,
(	31826	)	,
(	31117	)	,
(	30438	)	,
(	29789	)	,
(	29166	)	,
(	28569	)	,
(	27996	)	,
(	27445	)	,
(	26915	)	,
(	26406	)	,
(	25915	)	,
(	25442	)	,
(	24986	)	,
(	24546	)	,
(	24121	)	,
(	23711	)	,
(	23314	)	,
(	22930	)	,
(	22559	)	,
(	22199	)	,
(	21851	)	,
(	21513	)	,
(	21186	)	,
(	20868	)	,
(	20560	)	,
(	20261	)	,
(	19970	)	,
(	19687	)	,
(	19413	)	,
(	19145	)	,
(	18885	)	,
(	18632	)	,
(	18386	)	,
(	18146	)	,
(	17912	)	,
(	17684	)	,
(	17462	)	,
(	17245	)	,
(	17034	)	,
(	16827	)	,
(	16626	)	,
(	16429	)	,
(	16237	)	,
(	16049	)	,
(	15866	)	,
(	15687	)	,
(	15511	)	,
(	15340	)	,
(	15172	)	,
(	15008	)	,
(	14847	)	,
(	14690	)	,
(	14536	)	,
(	14385	)	,
(	14237	)	,
(	14093	)	,
(	13951	)	,
(	13812	)	,
(	13675	)	,
(	13542	)	,
(	13411	)	,
(	13282	)	,
(	13156	)	,
(	13032	)	,
(	12910	)	,
(	12791	)	,
(	12674	)	,
(	12559	)	,
(	12446	)	,
(	12335	)	,
(	12226	)	,
(	12119	)	,
(	12013	)	,
(	11910	)	,
(	11808	)	,
(	11708	)	,
(	11610	)	,
(	11513	)	,
(	11418	)	,
(	11324	)	,
(	11232	)	,
(	11142	)	,
(	11053	)	,
(	10965	)	,
(	10878	)	,
(	10793	)	,
(	10710	)	,
(	10627	)	,
(	10546	)	,
(	10466	)	,
(	10387	)	,
(	10309	)	,
(	10233	)	,
(	10158	)	,
(	10083	)	,
(	10010	)	,
(	9938	)	,
(	9867	)	,
(	9797	)	,
(	9727	)	,
(	9659	)	,
(	9592	)	,
(	9526	)	,
(	9460	)	,
(	9396	)	,
(	9332	)	,
(	9269	)	,
(	9207	)	,
(	9146	)	,
(	9085	)	,
(	9026	)	,
(	8967	)	,
(	8909	)	,
(	8852	)	,
(	8795	)	,
(	8739	)	,
(	8684	)	,
(	8629	)	,
(	8575	)	,
(	8522	)	,
(	8470	)	,
(	8418	)	,
(	8367	)	,
(	8316	)	,
(	8266	)	,
(	8216	)	,
(	8167	)	,
(	8119	)	,
(	8071	)	,
(	8024	)	,
(	7978	)	,
(	7931	)	,
(	7886	)	,
(	7841	)	,
(	7796	)	,
(	7752	)	,
(	7709	)	,
(	7665	)	,
(	7623	)	,
(	7581	)	,
(	7539	)	,
(	7498	)	,
(	7457	)	,
(	7416	)	,
(	7376	)	,
(	7337	)	,
(	7298	)	,
(	7259	)	,
(	7221	)	,
(	7183	)	,
(	7145	)	,
(	7108	)	,
(	7072	)	,
(	7035	)	,
(	6999	)	,
(	6964	)	,
(	6928	)	,
(	6893	)	,
(	6859	)	,
(	6824	)	,
(	6791	)	,
(	6757	)	,
(	6724	)	,
(	6691	)	,
(	6658	)	,
(	6626	)	,
(	6594	)	,
(	6562	)	,
(	6531	)	,
(	6500	)	,
(	6469	)	,
(	6438	)	,
(	6408	)	,
(	6378	)	,
(	6348	)	,
(	6319	)	,
(	6290	)	,
(	6261	)	,
(	6232	)	,
(	6204	)	,
(	6176	)	,
(	6148	)	,
(	6120	)	,
(	6093	)	,
(	6066	)	,
(	6039	)	,
(	6012	)	,
(	5986	)	,
(	5960	)	,
(	5934	)	,
(	5908	)	,
(	5882	)	,
(	5857	)	,
(	5832	)	,
(	5807	)	,
(	5782	)	,
(	5758	)	,
(	5734	)	,
(	5709	)	,
(	5686	)	,
(	5662	)	,
(	5638	)	,
(	5615	)	,
(	5592	)	,
(	5569	)	,
(	5546	)	,
(	5524	)	,
(	5501	)	,
(	5479	)	,
(	5457	)	,
(	5435	)	,
(	5414	)	,
(	5392	)	,
(	5371	)	,
(	5350	)	,
(	5329	)	,
(	5308	)	,
(	5287	)	,
(	5266	)	,
(	5246	)	,
(	5226	)	,
(	5206	)	,
(	5186	)	,
(	5166	)	,
(	5146	)	,
(	5127	)	,
(	5108	)	,
(	5088	)	,
(	5069	)	,
(	5050	)	,
(	5032	)	,
(	5013	)	,
(	4995	)	,
(	4976	)	,
(	4958	)	,
(	4940	)	,
(	4922	)	,
(	4904	)	,
(	4886	)	,
(	4869	)	,
(	4851	)	,
(	4834	)	,
(	4817	)	,
(	4799	)	,
(	4782	)	,
(	4766	)	,
(	4749	)	,
(	4732	)	,
(	4716	)	,
(	4699	)	,
(	4683	)	,
(	4667	)	,
(	4651	)	,
(	4635	)	,
(	4619	)	,
(	4603	)	,
(	4587	)	,
(	4572	)	,
(	4556	)	,
(	4541	)	,
(	4526	)	,
(	4511	)	,
(	4496	)	,
(	4481	)	,
(	4466	)	,
(	4451	)	,
(	4436	)	,
(	4422	)	,
(	4407	)	,
(	4393	)	,
(	4379	)	,
(	4364	)	,
(	4350	)	,
(	4336	)	,
(	4322	)	,
(	4309	)	,
(	4295	)	,
(	4281	)	,
(	4268	)	,
(	4254	)	,
(	4241	)	,
(	4227	)	,
(	4214	)	,
(	4201	)	,
(	4188	)	,
(	4175	)	,
(	4162	)	,
(	4149	)	,
(	4136	)	,
(	4123	)	,
(	4111	)	,
(	4098	)	,
(	4086	)	,
(	4073	)	,
(	4061	)	,
(	4049	)	,
(	4037	)	,
(	4025	)	,
(	4012	)	,
(	4000	)	,
(	3989	)	,
(	3977	)	,
(	3965	)	,
(	3953	)	,
(	3942	)	,
(	3930	)	,
(	3919	)	,
(	3907	)	,
(	3896	)	,
(	3884	)	,
(	3873	)	,
(	3862	)	,
(	3851	)	,
(	3840	)	,
(	3829	)	,
(	3818	)	,
(	3807	)	,
(	3796	)	,
(	3786	)	,
(	3775	)	,
(	3764	)	,
(	3754	)	,
(	3743	)	,
(	3733	)	,
(	3722	)	,
(	3712	)	,
(	3702	)	,
(	3691	)	,
(	3681	)	,
(	3671	)	,
(	3661	)	,
(	3651	)	,
(	3641	)	,
(	3631	)	,
(	3621	)	,
(	3612	)	,
(	3602	)	,
(	3592	)	,
(	3582	)	,
(	3573	)	,
(	3563	)	,
(	3554	)	,
(	3544	)	,
(	3535	)	,
(	3526	)	,
(	3516	)	,
(	3507	)	,
(	3498	)	,
(	3489	)	,
(	3480	)	,
(	3470	)	,
(	3461	)	,
(	3452	)	,
(	3444	)	,
(	3435	)	,
(	3426	)	,
(	3417	)	,
(	3408	)	,
(	3400	)	,
(	3391	)	,
(	3382	)	,
(	3374	)	,
(	3365	)	,
(	3357	)	,
(	3348	)	,
(	3340	)	,
(	3331	)	,
(	3323	)	,
(	3315	)	,
(	3306	)	,
(	3298	)	,
(	3290	)	,
(	3282	)	,
(	3274	)	,
(	3266	)	,
(	3258	)	,
(	3250	)	,
(	3242	)	,
(	3234	)	,
(	3226	)	,
(	3218	)	,
(	3210	)	,
(	3203	)	,
(	3195	)	,
(	3187	)	,
(	3180	)	,
(	3172	)	,
(	3164	)	,
(	3157	)	,
(	3149	)	,
(	3142	)	,
(	3134	)	,
(	3127	)	,
(	3120	)	,
(	3112	)	,
(	3105	)	,
(	3098	)	,
(	3091	)	,
(	3083	)	,
(	3076	)	,
(	3069	)	,
(	3062	)	,
(	3055	)	,
(	3048	)	,
(	3041	)	,
(	3034	)	,
(	3027	)	,
(	3020	)	,
(	3013	)	,
(	3006	)	,
(	2999	)	,
(	2993	)	,
(	2986	)	,
(	2979	)	,
(	2972	)	,
(	2966	)	,
(	2959	)	,
(	2952	)	,
(	2946	)	,
(	2939	)	,
(	2933	)	,
(	2926	)	,
(	2920	)	,
(	2913	)	,
(	2907	)	,
(	2900	)	,
(	2894	)	,
(	2888	)	,
(	2881	)	,
(	2875	)	,
(	2869	)	,
(	2863	)	,
(	2856	)	,
(	2850	)	,
(	2844	)	,
(	2838	)	,
(	2832	)	,
(	2826	)	,
(	2820	)	,
(	2814	)	,
(	2808	)	,
(	2802	)	,
(	2796	)	,
(	2790	)	,
(	2784	)	,
(	2778	)	,
(	2772	)	,
(	2766	)	,
(	2760	)	,
(	2755	)	,
(	2749	)	,
(	2743	)	,
(	2737	)	,
(	2732	)	,
(	2726	)	,
(	2720	)	,
(	2715	)	,
(	2709	)	,
(	2704	)	,
(	2698	)	,
(	2692	)	,
(	2687	)	,
(	2681	)	,
(	2676	)	,
(	2671	)	,
(	2665	)	,
(	2660	)	,
(	2654	)	,
(	2649	)	,
(	2644	)	,
(	2638	)	,
(	2633	)	,
(	2628	)	,
(	2622	)	,
(	2617	)	,
(	2612	)	,
(	2607	)	,
(	2602	)	,
(	2596	)	,
(	2591	)	,
(	2586	)	,
(	2581	)	,
(	2576	)	,
(	2571	)	,
(	2566	)	,
(	2561	)	,
(	2556	)	,
(	2551	)	,
(	2546	)	,
(	2541	)	,
(	2536	)	,
(	2531	)	,
(	2526	)	,
(	2521	)	,
(	2516	)	,
(	2511	)	,
(	2507	)	,
(	2502	)	,
(	2497	)	,
(	2492	)	,
(	2488	)	,
(	2483	)	,
(	2478	)	,
(	2473	)	,
(	2469	)	,
(	2464	)	,
(	2459	)	,
(	2455	)	,
(	2450	)	,
(	2446	)	,
(	2441	)	,
(	2436	)	,
(	2432	)	,
(	2427	)	,
(	2423	)	,
(	2418	)	,
(	2414	)	,
(	2409	)	,
(	2405	)	,
(	2400	)	,
(	2396	)	,
(	2392	)	,
(	2387	)	,
(	2383	)	,
(	2378	)	,
(	2374	)	,
(	2370	)	,
(	2365	)	,
(	2361	)	,
(	2357	)	,
(	2353	)	,
(	2348	)	,
(	2344	)	,
(	2340	)	,
(	2336	)	,
(	2331	)	,
(	2327	)	,
(	2323	)	,
(	2319	)	,
(	2315	)	,
(	2311	)	,
(	2307	)	,
(	2303	)	,
(	2298	)	,
(	2294	)	,
(	2290	)	,
(	2286	)	,
(	2282	)	,
(	2278	)	,
(	2274	)	,
(	2270	)	,
(	2266	)	,
(	2262	)	,
(	2258	)	,
(	2254	)	,
(	2250	)	,
(	2247	)	,
(	2243	)	,
(	2239	)	,
(	2235	)	,
(	2231	)	,
(	2227	)	,
(	2223	)	,
(	2220	)	,
(	2216	)	,
(	2212	)	,
(	2208	)	,
(	2204	)	,
(	2201	)	,
(	2197	)	,
(	2193	)	,
(	2189	)	,
(	2186	)	,
(	2182	)	,
(	2178	)	,
(	2175	)	,
(	2171	)	,
(	2167	)	,
(	2164	)	,
(	2160	)	,
(	2157	)	,
(	2153	)	,
(	2149	)	,
(	2146	)	,
(	2142	)	,
(	2139	)	,
(	2135	)	,
(	2132	)	,
(	2128	)	,
(	2125	)	,
(	2121	)	,
(	2118	)	,
(	2114	)	,
(	2111	)	,
(	2107	)	,
(	2104	)	,
(	2100	)	,
(	2097	)	,
(	2093	)	,
(	2090	)	,
(	2087	)	,
(	2083	)	,
(	2080	)	,
(	2077	)	,
(	2073	)	,
(	2070	)	,
(	2067	)	,
(	2063	)	,
(	2060	)	,
(	2057	)	,
(	2053	)	,
(	2050	)	,
(	2047	)	,
(	2043	)	,
(	2040	)	,
(	2037	)	,
(	2034	)	,
(	2031	)	,
(	2027	)	,
(	2024	)	,
(	2021	)	,
(	2018	)	,
(	2015	)	,
(	2011	)	,
(	2008	)	,
(	2005	)	,
(	2002	)	,
(	1999	)	,
(	1996	)	,
(	1993	)	,
(	1990	)	,
(	1986	)	,
(	1983	)	,
(	1980	)	,
(	1977	)	,
(	1974	)	,
(	1971	)	,
(	1968	)	,
(	1965	)	,
(	1962	)	,
(	1959	)	,
(	1956	)	,
(	1953	)	,
(	1950	)	,
(	1947	)	,
(	1944	)	,
(	1941	)	,
(	1938	)	,
(	1935	)	,
(	1932	)	,
(	1930	)	,
(	1927	)	,
(	1924	)	,
(	1921	)	,
(	1918	)	,
(	1915	)	,
(	1912	)	,
(	1909	)	,
(	1906	)	,
(	1904	)	,
(	1901	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1890	)	,
(	1887	)	,
(	1884	)	,
(	1881	)	,
(	1878	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1865	)	,
(	1862	)	,
(	1859	)	,
(	1856	)	,
(	1854	)	,
(	1851	)	,
(	1848	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1838	)	,
(	1835	)	,
(	1832	)	,
(	1830	)	,
(	1827	)	,
(	1824	)	,
(	1822	)	,
(	1819	)	,
(	1817	)	,
(	1814	)	,
(	1811	)	,
(	1809	)	,
(	1806	)	,
(	1804	)	,
(	1801	)	,
(	1799	)	,
(	1796	)	,
(	1794	)	,
(	1791	)	,
(	1788	)	,
(	1786	)	,
(	1783	)	,
(	1781	)	,
(	1778	)	,
(	1776	)	,
(	1773	)	,
(	1771	)	,
(	1768	)	,
(	1766	)	,
(	1764	)	,
(	1761	)	,
(	1759	)	,
(	1756	)	,
(	1754	)	,
(	1751	)	,
(	1749	)	,
(	1747	)	,
(	1744	)	,
(	1742	)	,
(	1739	)	,
(	1737	)	,
(	1735	)	,
(	1732	)	,
(	1730	)	,
(	1727	)	,
(	1725	)	,
(	1723	)	,
(	1720	)	,
(	1718	)	,
(	1716	)	,
(	1713	)	,
(	1711	)	,
(	1709	)	,
(	1706	)	,
(	1704	)	,
(	1702	)	,
(	1699	)	,
(	1697	)	,
(	1695	)	,
(	1693	)	,
(	1690	)	,
(	1688	)	,
(	1686	)	,
(	1684	)	,
(	1681	)	,
(	1679	)	,
(	1677	)	,
(	1675	)	,
(	1672	)	,
(	1670	)	,
(	1668	)	,
(	1666	)	,
(	1664	)	,
(	1661	)	,
(	1659	)	,
(	1657	)	,
(	1655	)	,
(	1653	)	,
(	1650	)	,
(	1648	)	,
(	1646	)	,
(	1644	)	,
(	1642	)	,
(	1640	)	,
(	1638	)	,
(	1635	)	,
(	1633	)	,
(	1631	)	,
(	1629	)	,
(	1627	)	,
(	1625	)	,
(	1623	)	,
(	1621	)	,
(	1619	)	,
(	1616	)	,
(	1614	)	,
(	1612	)	,
(	1610	)	,
(	1608	)	,
(	1606	)	,
(	1604	)	,
(	1602	)	,
(	1600	)	,
(	1598	)	,
(	1596	)	,
(	1594	)	,
(	1592	)	,
(	1590	)	,
(	1588	)	,
(	1586	)	,
(	1584	)	,
(	1582	)	,
(	1580	)	,
(	1578	)	,
(	1576	)	,
(	1574	)	,
(	1572	)	,
(	1570	)	,
(	1568	)	,
(	1566	)	,
(	1564	)	,
(	1562	)	,
(	1560	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1552	)	,
(	1550	)	,
(	1548	)	,
(	1547	)	,
(	1545	)	,
(	1543	)	,
(	1541	)	,
(	1539	)	,
(	1537	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1529	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1518	)	,
(	1516	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1507	)	,
(	1505	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1496	)	,
(	1495	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1486	)	,
(	1484	)	,
(	1482	)	,
(	1480	)	,
(	1479	)	,
(	1477	)	,
(	1475	)	,
(	1473	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1465	)	,
(	1463	)	,
(	1461	)	,
(	1459	)	,
(	1458	)	,
(	1456	)	,
(	1454	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1447	)	,
(	1446	)	,
(	1444	)	,
(	1442	)	,
(	1441	)	,
(	1439	)	,
(	1437	)	,
(	1436	)	,
(	1434	)	,
(	1432	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1426	)	,
(	1424	)	,
(	1422	)	,
(	1421	)	,
(	1419	)	,
(	1418	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1408	)	,
(	1406	)	,
(	1405	)	,
(	1403	)	,
(	1401	)	,
(	1400	)	,
(	1398	)	,
(	1397	)	,
(	1395	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1389	)	,
(	1387	)	,
(	1386	)	,
(	1384	)	,
(	1383	)	,
(	1381	)	,
(	1380	)	,
(	1378	)	,
(	1376	)	,
(	1375	)	,
(	1373	)	,
(	1372	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1364	)	,
(	1363	)	,
(	1361	)	,
(	1360	)	,
(	1358	)	,
(	1357	)	,
(	1355	)	,
(	1354	)	,
(	1352	)	,
(	1351	)	,
(	1349	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1337	)	,
(	1336	)	,
(	1335	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1323	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1306	)	,
(	1305	)	,
(	1303	)	,
(	1302	)	,
(	1300	)	,
(	1299	)	,
(	1298	)	,
(	1296	)	,
(	1295	)	,
(	1294	)	,
(	1292	)	,
(	1291	)	,
(	1289	)	,
(	1288	)	,
(	1287	)	,
(	1285	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1272	)	,
(	1271	)	,
(	1269	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1252	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1246	)	,
(	1245	)	,
(	1243	)	,
(	1242	)	,
(	1241	)	,
(	1240	)	,
(	1238	)	,
(	1237	)	,
(	1236	)	,
(	1235	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1230	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1220	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1215	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1203	)	,
(	1201	)	,
(	1200	)	,
(	1199	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1188	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1183	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1167	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1162	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1146	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1141	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1135	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1115	)	,
(	1114	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	938	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	929	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	399	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	398	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	397	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	396	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	395	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	394	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	393	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	392	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	391	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	390	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	389	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	388	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	387	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	386	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	385	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	384	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	383	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	382	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	381	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	380	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	379	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	378	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	377	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	376	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	375	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	374	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	373	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	372	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	371	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	370	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	369	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	368	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	367	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	366	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	365	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	364	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	363	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	
			


);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));
	
	
	process(voltage)
	begin
		if(unsigned(voltage) <= 414) then
			err_flag <= '1';
		else
			err_flag <= '0';
		end if;
	end process;

end behavior;
