LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2frequency IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      frequency      :  OUT   natural
		);		
END voltage2frequency;

ARCHITECTURE behavior OF voltage2frequency IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2f_LUT : array_1d := (

(	3333	)	,
(	3335	)	,
(	3337	)	,
(	3338	)	,
(	3340	)	,
(	3341	)	,
(	3343	)	,
(	3345	)	,
(	3346	)	,
(	3348	)	,
(	3350	)	,
(	3351	)	,
(	3353	)	,
(	3354	)	,
(	3356	)	,
(	3358	)	,
(	3359	)	,
(	3361	)	,
(	3362	)	,
(	3364	)	,
(	3366	)	,
(	3367	)	,
(	3369	)	,
(	3371	)	,
(	3372	)	,
(	3374	)	,
(	3375	)	,
(	3377	)	,
(	3379	)	,
(	3380	)	,
(	3382	)	,
(	3384	)	,
(	3385	)	,
(	3387	)	,
(	3388	)	,
(	3390	)	,
(	3392	)	,
(	3393	)	,
(	3395	)	,
(	3397	)	,
(	3398	)	,
(	3400	)	,
(	3401	)	,
(	3403	)	,
(	3405	)	,
(	3406	)	,
(	3408	)	,
(	3409	)	,
(	3411	)	,
(	3413	)	,
(	3414	)	,
(	3416	)	,
(	3418	)	,
(	3419	)	,
(	3421	)	,
(	3422	)	,
(	3424	)	,
(	3426	)	,
(	3427	)	,
(	3429	)	,
(	3431	)	,
(	3432	)	,
(	3434	)	,
(	3435	)	,
(	3437	)	,
(	3439	)	,
(	3440	)	,
(	3442	)	,
(	3443	)	,
(	3445	)	,
(	3447	)	,
(	3448	)	,
(	3450	)	,
(	3452	)	,
(	3453	)	,
(	3455	)	,
(	3456	)	,
(	3458	)	,
(	3460	)	,
(	3461	)	,
(	3463	)	,
(	3465	)	,
(	3466	)	,
(	3468	)	,
(	3469	)	,
(	3471	)	,
(	3473	)	,
(	3474	)	,
(	3476	)	,
(	3478	)	,
(	3479	)	,
(	3481	)	,
(	3482	)	,
(	3484	)	,
(	3486	)	,
(	3487	)	,
(	3489	)	,
(	3490	)	,
(	3492	)	,
(	3494	)	,
(	3495	)	,
(	3497	)	,
(	3499	)	,
(	3500	)	,
(	3502	)	,
(	3503	)	,
(	3505	)	,
(	3507	)	,
(	3508	)	,
(	3510	)	,
(	3512	)	,
(	3513	)	,
(	3515	)	,
(	3516	)	,
(	3518	)	,
(	3520	)	,
(	3521	)	,
(	3523	)	,
(	3524	)	,
(	3526	)	,
(	3528	)	,
(	3529	)	,
(	3531	)	,
(	3533	)	,
(	3534	)	,
(	3536	)	,
(	3537	)	,
(	3539	)	,
(	3541	)	,
(	3542	)	,
(	3544	)	,
(	3546	)	,
(	3547	)	,
(	3549	)	,
(	3550	)	,
(	3552	)	,
(	3554	)	,
(	3555	)	,
(	3557	)	,
(	3559	)	,
(	3560	)	,
(	3562	)	,
(	3563	)	,
(	3565	)	,
(	3567	)	,
(	3568	)	,
(	3570	)	,
(	3571	)	,
(	3573	)	,
(	3575	)	,
(	3576	)	,
(	3578	)	,
(	3580	)	,
(	3581	)	,
(	3583	)	,
(	3584	)	,
(	3586	)	,
(	3588	)	,
(	3589	)	,
(	3591	)	,
(	3593	)	,
(	3594	)	,
(	3596	)	,
(	3597	)	,
(	3599	)	,
(	3601	)	,
(	3602	)	,
(	3604	)	,
(	3605	)	,
(	3607	)	,
(	3609	)	,
(	3610	)	,
(	3612	)	,
(	3614	)	,
(	3615	)	,
(	3617	)	,
(	3618	)	,
(	3620	)	,
(	3622	)	,
(	3623	)	,
(	3625	)	,
(	3627	)	,
(	3628	)	,
(	3630	)	,
(	3631	)	,
(	3633	)	,
(	3635	)	,
(	3636	)	,
(	3638	)	,
(	3640	)	,
(	3641	)	,
(	3643	)	,
(	3644	)	,
(	3646	)	,
(	3648	)	,
(	3649	)	,
(	3651	)	,
(	3652	)	,
(	3654	)	,
(	3656	)	,
(	3657	)	,
(	3659	)	,
(	3661	)	,
(	3662	)	,
(	3664	)	,
(	3665	)	,
(	3667	)	,
(	3669	)	,
(	3670	)	,
(	3672	)	,
(	3674	)	,
(	3675	)	,
(	3677	)	,
(	3678	)	,
(	3680	)	,
(	3682	)	,
(	3683	)	,
(	3685	)	,
(	3686	)	,
(	3688	)	,
(	3690	)	,
(	3691	)	,
(	3693	)	,
(	3695	)	,
(	3696	)	,
(	3698	)	,
(	3699	)	,
(	3701	)	,
(	3703	)	,
(	3704	)	,
(	3706	)	,
(	3708	)	,
(	3709	)	,
(	3711	)	,
(	3712	)	,
(	3714	)	,
(	3716	)	,
(	3717	)	,
(	3719	)	,
(	3721	)	,
(	3722	)	,
(	3724	)	,
(	3725	)	,
(	3727	)	,
(	3729	)	,
(	3730	)	,
(	3732	)	,
(	3733	)	,
(	3735	)	,
(	3737	)	,
(	3738	)	,
(	3740	)	,
(	3742	)	,
(	3743	)	,
(	3745	)	,
(	3746	)	,
(	3748	)	,
(	3750	)	,
(	3751	)	,
(	3753	)	,
(	3755	)	,
(	3756	)	,
(	3758	)	,
(	3759	)	,
(	3761	)	,
(	3763	)	,
(	3764	)	,
(	3766	)	,
(	3767	)	,
(	3769	)	,
(	3771	)	,
(	3772	)	,
(	3774	)	,
(	3776	)	,
(	3777	)	,
(	3779	)	,
(	3780	)	,
(	3782	)	,
(	3784	)	,
(	3785	)	,
(	3787	)	,
(	3789	)	,
(	3790	)	,
(	3792	)	,
(	3793	)	,
(	3795	)	,
(	3797	)	,
(	3798	)	,
(	3800	)	,
(	3802	)	,
(	3803	)	,
(	3805	)	,
(	3806	)	,
(	3808	)	,
(	3810	)	,
(	3811	)	,
(	3813	)	,
(	3814	)	,
(	3816	)	,
(	3818	)	,
(	3819	)	,
(	3821	)	,
(	3823	)	,
(	3824	)	,
(	3826	)	,
(	3827	)	,
(	3829	)	,
(	3831	)	,
(	3832	)	,
(	3834	)	,
(	3836	)	,
(	3837	)	,
(	3839	)	,
(	3840	)	,
(	3842	)	,
(	3844	)	,
(	3845	)	,
(	3847	)	,
(	3848	)	,
(	3850	)	,
(	3852	)	,
(	3853	)	,
(	3855	)	,
(	3857	)	,
(	3858	)	,
(	3860	)	,
(	3861	)	,
(	3863	)	,
(	3865	)	,
(	3866	)	,
(	3868	)	,
(	3870	)	,
(	3871	)	,
(	3873	)	,
(	3874	)	,
(	3876	)	,
(	3878	)	,
(	3879	)	,
(	3881	)	,
(	3883	)	,
(	3884	)	,
(	3886	)	,
(	3887	)	,
(	3889	)	,
(	3891	)	,
(	3892	)	,
(	3894	)	,
(	3895	)	,
(	3897	)	,
(	3899	)	,
(	3900	)	,
(	3902	)	,
(	3904	)	,
(	3905	)	,
(	3907	)	,
(	3908	)	,
(	3910	)	,
(	3912	)	,
(	3913	)	,
(	3915	)	,
(	3917	)	,
(	3918	)	,
(	3920	)	,
(	3921	)	,
(	3923	)	,
(	3925	)	,
(	3926	)	,
(	3928	)	,
(	3929	)	,
(	3931	)	,
(	3933	)	,
(	3934	)	,
(	3936	)	,
(	3938	)	,
(	3939	)	,
(	3941	)	,
(	3942	)	,
(	3944	)	,
(	3946	)	,
(	3947	)	,
(	3949	)	,
(	3951	)	,
(	3952	)	,
(	3954	)	,
(	3955	)	,
(	3957	)	,
(	3959	)	,
(	3960	)	,
(	3962	)	,
(	3964	)	,
(	3965	)	,
(	3967	)	,
(	3968	)	,
(	3970	)	,
(	3972	)	,
(	3973	)	,
(	3975	)	,
(	3976	)	,
(	3978	)	,
(	3980	)	,
(	3981	)	,
(	3983	)	,
(	3985	)	,
(	3986	)	,
(	3988	)	,
(	3989	)	,
(	3991	)	,
(	3993	)	,
(	3994	)	,
(	3996	)	,
(	3998	)	,
(	3999	)	,
(	4001	)	,
(	4002	)	,
(	4004	)	,
(	4006	)	,
(	4007	)	,
(	4009	)	,
(	4010	)	,
(	4012	)	,
(	4014	)	,
(	4015	)	,
(	4017	)	,
(	4019	)	,
(	4020	)	,
(	4022	)	,
(	4023	)	,
(	4025	)	,
(	4027	)	,
(	4028	)	,
(	4030	)	,
(	4032	)	,
(	4033	)	,
(	4035	)	,
(	4036	)	,
(	4038	)	,
(	4040	)	,
(	4041	)	,
(	4043	)	,
(	4045	)	,
(	4046	)	,
(	4048	)	,
(	4049	)	,
(	4051	)	,
(	4053	)	,
(	4054	)	,
(	4056	)	,
(	4057	)	,
(	4059	)	,
(	4061	)	,
(	4062	)	,
(	4064	)	,
(	4066	)	,
(	4067	)	,
(	4069	)	,
(	4070	)	,
(	4072	)	,
(	4074	)	,
(	4075	)	,
(	4077	)	,
(	4079	)	,
(	4080	)	,
(	4082	)	,
(	4083	)	,
(	4085	)	,
(	4087	)	,
(	4088	)	,
(	4090	)	,
(	4091	)	,
(	4093	)	,
(	4095	)	,
(	4096	)	,
(	4098	)	,
(	4100	)	,
(	4101	)	,
(	4103	)	,
(	4104	)	,
(	4106	)	,
(	4108	)	,
(	4109	)	,
(	4111	)	,
(	4113	)	,
(	4114	)	,
(	4116	)	,
(	4117	)	,
(	4119	)	,
(	4121	)	,
(	4122	)	,
(	4124	)	,
(	4126	)	,
(	4127	)	,
(	4129	)	,
(	4130	)	,
(	4132	)	,
(	4134	)	,
(	4135	)	,
(	4137	)	,
(	4138	)	,
(	4140	)	,
(	4142	)	,
(	4143	)	,
(	4145	)	,
(	4147	)	,
(	4148	)	,
(	4150	)	,
(	4151	)	,
(	4153	)	,
(	4155	)	,
(	4156	)	,
(	4158	)	,
(	4160	)	,
(	4161	)	,
(	4163	)	,
(	4164	)	,
(	4166	)	,
(	4168	)	,
(	4169	)	,
(	4171	)	,
(	4172	)	,
(	4174	)	,
(	4176	)	,
(	4177	)	,
(	4179	)	,
(	4181	)	,
(	4182	)	,
(	4184	)	,
(	4185	)	,
(	4187	)	,
(	4189	)	,
(	4190	)	,
(	4192	)	,
(	4194	)	,
(	4195	)	,
(	4197	)	,
(	4198	)	,
(	4200	)	,
(	4202	)	,
(	4203	)	,
(	4205	)	,
(	4207	)	,
(	4208	)	,
(	4210	)	,
(	4211	)	,
(	4213	)	,
(	4215	)	,
(	4216	)	,
(	4218	)	,
(	4219	)	,
(	4221	)	,
(	4223	)	,
(	4224	)	,
(	4226	)	,
(	4228	)	,
(	4229	)	,
(	4231	)	,
(	4232	)	,
(	4234	)	,
(	4236	)	,
(	4237	)	,
(	4239	)	,
(	4241	)	,
(	4242	)	,
(	4244	)	,
(	4245	)	,
(	4247	)	,
(	4249	)	,
(	4250	)	,
(	4252	)	,
(	4253	)	,
(	4255	)	,
(	4257	)	,
(	4258	)	,
(	4260	)	,
(	4262	)	,
(	4263	)	,
(	4265	)	,
(	4266	)	,
(	4268	)	,
(	4270	)	,
(	4271	)	,
(	4273	)	,
(	4275	)	,
(	4276	)	,
(	4278	)	,
(	4279	)	,
(	4281	)	,
(	4283	)	,
(	4284	)	,
(	4286	)	,
(	4288	)	,
(	4289	)	,
(	4291	)	,
(	4292	)	,
(	4294	)	,
(	4296	)	,
(	4297	)	,
(	4299	)	,
(	4300	)	,
(	4302	)	,
(	4304	)	,
(	4305	)	,
(	4307	)	,
(	4309	)	,
(	4310	)	,
(	4312	)	,
(	4313	)	,
(	4315	)	,
(	4317	)	,
(	4318	)	,
(	4320	)	,
(	4322	)	,
(	4323	)	,
(	4325	)	,
(	4326	)	,
(	4328	)	,
(	4330	)	,
(	4331	)	,
(	4333	)	,
(	4334	)	,
(	4336	)	,
(	4338	)	,
(	4339	)	,
(	4341	)	,
(	4343	)	,
(	4344	)	,
(	4346	)	,
(	4347	)	,
(	4349	)	,
(	4351	)	,
(	4352	)	,
(	4354	)	,
(	4356	)	,
(	4357	)	,
(	4359	)	,
(	4360	)	,
(	4362	)	,
(	4364	)	,
(	4365	)	,
(	4367	)	,
(	4369	)	,
(	4370	)	,
(	4372	)	,
(	4373	)	,
(	4375	)	,
(	4377	)	,
(	4378	)	,
(	4380	)	,
(	4381	)	,
(	4383	)	,
(	4385	)	,
(	4386	)	,
(	4388	)	,
(	4390	)	,
(	4391	)	,
(	4393	)	,
(	4394	)	,
(	4396	)	,
(	4398	)	,
(	4399	)	,
(	4401	)	,
(	4403	)	,
(	4404	)	,
(	4406	)	,
(	4407	)	,
(	4409	)	,
(	4411	)	,
(	4412	)	,
(	4414	)	,
(	4415	)	,
(	4417	)	,
(	4419	)	,
(	4420	)	,
(	4422	)	,
(	4424	)	,
(	4425	)	,
(	4427	)	,
(	4428	)	,
(	4430	)	,
(	4432	)	,
(	4433	)	,
(	4435	)	,
(	4437	)	,
(	4438	)	,
(	4440	)	,
(	4441	)	,
(	4443	)	,
(	4445	)	,
(	4446	)	,
(	4448	)	,
(	4450	)	,
(	4451	)	,
(	4453	)	,
(	4454	)	,
(	4456	)	,
(	4458	)	,
(	4459	)	,
(	4461	)	,
(	4462	)	,
(	4464	)	,
(	4466	)	,
(	4467	)	,
(	4469	)	,
(	4471	)	,
(	4472	)	,
(	4474	)	,
(	4475	)	,
(	4477	)	,
(	4479	)	,
(	4480	)	,
(	4482	)	,
(	4484	)	,
(	4485	)	,
(	4487	)	,
(	4488	)	,
(	4490	)	,
(	4492	)	,
(	4493	)	,
(	4495	)	,
(	4496	)	,
(	4498	)	,
(	4500	)	,
(	4501	)	,
(	4503	)	,
(	4505	)	,
(	4506	)	,
(	4508	)	,
(	4509	)	,
(	4511	)	,
(	4513	)	,
(	4514	)	,
(	4516	)	,
(	4518	)	,
(	4519	)	,
(	4521	)	,
(	4522	)	,
(	4524	)	,
(	4526	)	,
(	4527	)	,
(	4529	)	,
(	4531	)	,
(	4532	)	,
(	4534	)	,
(	4535	)	,
(	4537	)	,
(	4539	)	,
(	4540	)	,
(	4542	)	,
(	4543	)	,
(	4545	)	,
(	4547	)	,
(	4548	)	,
(	4550	)	,
(	4552	)	,
(	4553	)	,
(	4555	)	,
(	4556	)	,
(	4558	)	,
(	4560	)	,
(	4561	)	,
(	4563	)	,
(	4565	)	,
(	4566	)	,
(	4568	)	,
(	4569	)	,
(	4571	)	,
(	4573	)	,
(	4574	)	,
(	4576	)	,
(	4577	)	,
(	4579	)	,
(	4581	)	,
(	4582	)	,
(	4584	)	,
(	4586	)	,
(	4587	)	,
(	4589	)	,
(	4590	)	,
(	4592	)	,
(	4594	)	,
(	4595	)	,
(	4597	)	,
(	4599	)	,
(	4600	)	,
(	4602	)	,
(	4603	)	,
(	4605	)	,
(	4607	)	,
(	4608	)	,
(	4610	)	,
(	4612	)	,
(	4613	)	,
(	4615	)	,
(	4616	)	,
(	4618	)	,
(	4620	)	,
(	4621	)	,
(	4623	)	,
(	4624	)	,
(	4626	)	,
(	4628	)	,
(	4629	)	,
(	4631	)	,
(	4633	)	,
(	4634	)	,
(	4636	)	,
(	4637	)	,
(	4639	)	,
(	4641	)	,
(	4642	)	,
(	4644	)	,
(	4646	)	,
(	4647	)	,
(	4649	)	,
(	4650	)	,
(	4652	)	,
(	4654	)	,
(	4655	)	,
(	4657	)	,
(	4658	)	,
(	4660	)	,
(	4662	)	,
(	4663	)	,
(	4665	)	,
(	4667	)	,
(	4668	)	,
(	4670	)	,
(	4671	)	,
(	4673	)	,
(	4675	)	,
(	4676	)	,
(	4678	)	,
(	4680	)	,
(	4681	)	,
(	4683	)	,
(	4684	)	,
(	4686	)	,
(	4688	)	,
(	4689	)	,
(	4691	)	,
(	4693	)	,
(	4694	)	,
(	4696	)	,
(	4697	)	,
(	4699	)	,
(	4701	)	,
(	4702	)	,
(	4704	)	,
(	4705	)	,
(	4707	)	,
(	4709	)	,
(	4710	)	,
(	4712	)	,
(	4714	)	,
(	4715	)	,
(	4717	)	,
(	4718	)	,
(	4720	)	,
(	4722	)	,
(	4723	)	,
(	4725	)	,
(	4727	)	,
(	4728	)	,
(	4730	)	,
(	4731	)	,
(	4733	)	,
(	4735	)	,
(	4736	)	,
(	4738	)	,
(	4739	)	,
(	4741	)	,
(	4743	)	,
(	4744	)	,
(	4746	)	,
(	4748	)	,
(	4749	)	,
(	4751	)	,
(	4752	)	,
(	4754	)	,
(	4756	)	,
(	4757	)	,
(	4759	)	,
(	4761	)	,
(	4762	)	,
(	4764	)	,
(	4765	)	,
(	4767	)	,
(	4769	)	,
(	4770	)	,
(	4772	)	,
(	4774	)	,
(	4775	)	,
(	4777	)	,
(	4778	)	,
(	4780	)	,
(	4782	)	,
(	4783	)	,
(	4785	)	,
(	4786	)	,
(	4788	)	,
(	4790	)	,
(	4791	)	,
(	4793	)	,
(	4795	)	,
(	4796	)	,
(	4798	)	,
(	4799	)	,
(	4801	)	,
(	4803	)	,
(	4804	)	,
(	4806	)	,
(	4808	)	,
(	4809	)	,
(	4811	)	,
(	4812	)	,
(	4814	)	,
(	4816	)	,
(	4817	)	,
(	4819	)	,
(	4820	)	,
(	4822	)	,
(	4824	)	,
(	4825	)	,
(	4827	)	,
(	4829	)	,
(	4830	)	,
(	4832	)	,
(	4833	)	,
(	4835	)	,
(	4837	)	,
(	4838	)	,
(	4840	)	,
(	4842	)	,
(	4843	)	,
(	4845	)	,
(	4846	)	,
(	4848	)	,
(	4850	)	,
(	4851	)	,
(	4853	)	,
(	4855	)	,
(	4856	)	,
(	4858	)	,
(	4859	)	,
(	4861	)	,
(	4863	)	,
(	4864	)	,
(	4866	)	,
(	4867	)	,
(	4869	)	,
(	4871	)	,
(	4872	)	,
(	4874	)	,
(	4876	)	,
(	4877	)	,
(	4879	)	,
(	4880	)	,
(	4882	)	,
(	4884	)	,
(	4885	)	,
(	4887	)	,
(	4889	)	,
(	4890	)	,
(	4892	)	,
(	4893	)	,
(	4895	)	,
(	4897	)	,
(	4898	)	,
(	4900	)	,
(	4901	)	,
(	4903	)	,
(	4905	)	,
(	4906	)	,
(	4908	)	,
(	4910	)	,
(	4911	)	,
(	4913	)	,
(	4914	)	,
(	4916	)	,
(	4918	)	,
(	4919	)	,
(	4921	)	,
(	4923	)	,
(	4924	)	,
(	4926	)	,
(	4927	)	,
(	4929	)	,
(	4931	)	,
(	4932	)	,
(	4934	)	,
(	4936	)	,
(	4937	)	,
(	4939	)	,
(	4940	)	,
(	4942	)	,
(	4944	)	,
(	4945	)	,
(	4947	)	,
(	4948	)	,
(	4950	)	,
(	4952	)	,
(	4953	)	,
(	4955	)	,
(	4957	)	,
(	4958	)	,
(	4960	)	,
(	4961	)	,
(	4963	)	,
(	4965	)	,
(	4966	)	,
(	4968	)	,
(	4970	)	,
(	4971	)	,
(	4973	)	,
(	4974	)	,
(	4976	)	,
(	4978	)	,
(	4979	)	,
(	4981	)	,
(	4982	)	,
(	4984	)	,
(	4986	)	,
(	4987	)	,
(	4989	)	,
(	4991	)	,
(	4992	)	,
(	4994	)	,
(	4995	)	,
(	4997	)	,
(	4999	)	,
(	5000	)	,
(	5002	)	,
(	5004	)	,
(	5005	)	,
(	5007	)	,
(	5008	)	,
(	5010	)	,
(	5012	)	,
(	5013	)	,
(	5015	)	,
(	5017	)	,
(	5018	)	,
(	5020	)	,
(	5021	)	,
(	5023	)	,
(	5025	)	,
(	5026	)	,
(	5028	)	,
(	5029	)	,
(	5031	)	,
(	5033	)	,
(	5034	)	,
(	5036	)	,
(	5038	)	,
(	5039	)	,
(	5041	)	,
(	5042	)	,
(	5044	)	,
(	5046	)	,
(	5047	)	,
(	5049	)	,
(	5051	)	,
(	5052	)	,
(	5054	)	,
(	5055	)	,
(	5057	)	,
(	5059	)	,
(	5060	)	,
(	5062	)	,
(	5063	)	,
(	5065	)	,
(	5067	)	,
(	5068	)	,
(	5070	)	,
(	5072	)	,
(	5073	)	,
(	5075	)	,
(	5076	)	,
(	5078	)	,
(	5080	)	,
(	5081	)	,
(	5083	)	,
(	5085	)	,
(	5086	)	,
(	5088	)	,
(	5089	)	,
(	5091	)	,
(	5093	)	,
(	5094	)	,
(	5096	)	,
(	5098	)	,
(	5099	)	,
(	5101	)	,
(	5102	)	,
(	5104	)	,
(	5106	)	,
(	5107	)	,
(	5109	)	,
(	5110	)	,
(	5112	)	,
(	5114	)	,
(	5115	)	,
(	5117	)	,
(	5119	)	,
(	5120	)	,
(	5122	)	,
(	5123	)	,
(	5125	)	,
(	5127	)	,
(	5128	)	,
(	5130	)	,
(	5132	)	,
(	5133	)	,
(	5135	)	,
(	5136	)	,
(	5138	)	,
(	5140	)	,
(	5141	)	,
(	5143	)	,
(	5144	)	,
(	5146	)	,
(	5148	)	,
(	5149	)	,
(	5151	)	,
(	5153	)	,
(	5154	)	,
(	5156	)	,
(	5157	)	,
(	5159	)	,
(	5161	)	,
(	5162	)	,
(	5164	)	,
(	5166	)	,
(	5167	)	,
(	5169	)	,
(	5170	)	,
(	5172	)	,
(	5174	)	,
(	5175	)	,
(	5177	)	,
(	5179	)	,
(	5180	)	,
(	5182	)	,
(	5183	)	,
(	5185	)	,
(	5187	)	,
(	5188	)	,
(	5190	)	,
(	5191	)	,
(	5193	)	,
(	5195	)	,
(	5196	)	,
(	5198	)	,
(	5200	)	,
(	5201	)	,
(	5203	)	,
(	5204	)	,
(	5206	)	,
(	5208	)	,
(	5209	)	,
(	5211	)	,
(	5213	)	,
(	5214	)	,
(	5216	)	,
(	5217	)	,
(	5219	)	,
(	5221	)	,
(	5222	)	,
(	5224	)	,
(	5225	)	,
(	5227	)	,
(	5229	)	,
(	5230	)	,
(	5232	)	,
(	5234	)	,
(	5235	)	,
(	5237	)	,
(	5238	)	,
(	5240	)	,
(	5242	)	,
(	5243	)	,
(	5245	)	,
(	5247	)	,
(	5248	)	,
(	5250	)	,
(	5251	)	,
(	5253	)	,
(	5255	)	,
(	5256	)	,
(	5258	)	,
(	5260	)	,
(	5261	)	,
(	5263	)	,
(	5264	)	,
(	5266	)	,
(	5268	)	,
(	5269	)	,
(	5271	)	,
(	5272	)	,
(	5274	)	,
(	5276	)	,
(	5277	)	,
(	5279	)	,
(	5281	)	,
(	5282	)	,
(	5284	)	,
(	5285	)	,
(	5287	)	,
(	5289	)	,
(	5290	)	,
(	5292	)	,
(	5294	)	,
(	5295	)	,
(	5297	)	,
(	5298	)	,
(	5300	)	,
(	5302	)	,
(	5303	)	,
(	5305	)	,
(	5306	)	,
(	5308	)	,
(	5310	)	,
(	5311	)	,
(	5313	)	,
(	5315	)	,
(	5316	)	,
(	5318	)	,
(	5319	)	,
(	5321	)	,
(	5323	)	,
(	5324	)	,
(	5326	)	,
(	5328	)	,
(	5329	)	,
(	5331	)	,
(	5332	)	,
(	5334	)	,
(	5336	)	,
(	5337	)	,
(	5339	)	,
(	5341	)	,
(	5342	)	,
(	5344	)	,
(	5345	)	,
(	5347	)	,
(	5349	)	,
(	5350	)	,
(	5352	)	,
(	5353	)	,
(	5355	)	,
(	5357	)	,
(	5358	)	,
(	5360	)	,
(	5362	)	,
(	5363	)	,
(	5365	)	,
(	5366	)	,
(	5368	)	,
(	5370	)	,
(	5371	)	,
(	5373	)	,
(	5375	)	,
(	5376	)	,
(	5378	)	,
(	5379	)	,
(	5381	)	,
(	5383	)	,
(	5384	)	,
(	5386	)	,
(	5387	)	,
(	5389	)	,
(	5391	)	,
(	5392	)	,
(	5394	)	,
(	5396	)	,
(	5397	)	,
(	5399	)	,
(	5400	)	,
(	5402	)	,
(	5404	)	,
(	5405	)	,
(	5407	)	,
(	5409	)	,
(	5410	)	,
(	5412	)	,
(	5413	)	,
(	5415	)	,
(	5417	)	,
(	5418	)	,
(	5420	)	,
(	5422	)	,
(	5423	)	,
(	5425	)	,
(	5426	)	,
(	5428	)	,
(	5430	)	,
(	5431	)	,
(	5433	)	,
(	5434	)	,
(	5436	)	,
(	5438	)	,
(	5439	)	,
(	5441	)	,
(	5443	)	,
(	5444	)	,
(	5446	)	,
(	5447	)	,
(	5449	)	,
(	5451	)	,
(	5452	)	,
(	5454	)	,
(	5456	)	,
(	5457	)	,
(	5459	)	,
(	5460	)	,
(	5462	)	,
(	5464	)	,
(	5465	)	,
(	5467	)	,
(	5468	)	,
(	5470	)	,
(	5472	)	,
(	5473	)	,
(	5475	)	,
(	5477	)	,
(	5478	)	,
(	5480	)	,
(	5481	)	,
(	5483	)	,
(	5485	)	,
(	5486	)	,
(	5488	)	,
(	5490	)	,
(	5491	)	,
(	5493	)	,
(	5494	)	,
(	5496	)	,
(	5498	)	,
(	5499	)	,
(	5501	)	,
(	5503	)	,
(	5504	)	,
(	5506	)	,
(	5507	)	,
(	5509	)	,
(	5511	)	,
(	5512	)	,
(	5514	)	,
(	5515	)	,
(	5517	)	,
(	5519	)	,
(	5520	)	,
(	5522	)	,
(	5524	)	,
(	5525	)	,
(	5527	)	,
(	5528	)	,
(	5530	)	,
(	5532	)	,
(	5533	)	,
(	5535	)	,
(	5537	)	,
(	5538	)	,
(	5540	)	,
(	5541	)	,
(	5543	)	,
(	5545	)	,
(	5546	)	,
(	5548	)	,
(	5549	)	,
(	5551	)	,
(	5553	)	,
(	5554	)	,
(	5556	)	,
(	5558	)	,
(	5559	)	,
(	5561	)	,
(	5562	)	,
(	5564	)	,
(	5566	)	,
(	5567	)	,
(	5569	)	,
(	5571	)	,
(	5572	)	,
(	5574	)	,
(	5575	)	,
(	5577	)	,
(	5579	)	,
(	5580	)	,
(	5582	)	,
(	5584	)	,
(	5585	)	,
(	5587	)	,
(	5588	)	,
(	5590	)	,
(	5592	)	,
(	5593	)	,
(	5595	)	,
(	5596	)	,
(	5598	)	,
(	5600	)	,
(	5601	)	,
(	5603	)	,
(	5605	)	,
(	5606	)	,
(	5608	)	,
(	5609	)	,
(	5611	)	,
(	5613	)	,
(	5614	)	,
(	5616	)	,
(	5618	)	,
(	5619	)	,
(	5621	)	,
(	5622	)	,
(	5624	)	,
(	5626	)	,
(	5627	)	,
(	5629	)	,
(	5630	)	,
(	5632	)	,
(	5634	)	,
(	5635	)	,
(	5637	)	,
(	5639	)	,
(	5640	)	,
(	5642	)	,
(	5643	)	,
(	5645	)	,
(	5647	)	,
(	5648	)	,
(	5650	)	,
(	5652	)	,
(	5653	)	,
(	5655	)	,
(	5656	)	,
(	5658	)	,
(	5660	)	,
(	5661	)	,
(	5663	)	,
(	5665	)	,
(	5666	)	,
(	5668	)	,
(	5669	)	,
(	5671	)	,
(	5673	)	,
(	5674	)	,
(	5676	)	,
(	5677	)	,
(	5679	)	,
(	5681	)	,
(	5682	)	,
(	5684	)	,
(	5686	)	,
(	5687	)	,
(	5689	)	,
(	5690	)	,
(	5692	)	,
(	5694	)	,
(	5695	)	,
(	5697	)	,
(	5699	)	,
(	5700	)	,
(	5702	)	,
(	5703	)	,
(	5705	)	,
(	5707	)	,
(	5708	)	,
(	5710	)	,
(	5711	)	,
(	5713	)	,
(	5715	)	,
(	5716	)	,
(	5718	)	,
(	5720	)	,
(	5721	)	,
(	5723	)	,
(	5724	)	,
(	5726	)	,
(	5728	)	,
(	5729	)	,
(	5731	)	,
(	5733	)	,
(	5734	)	,
(	5736	)	,
(	5737	)	,
(	5739	)	,
(	5741	)	,
(	5742	)	,
(	5744	)	,
(	5746	)	,
(	5747	)	,
(	5749	)	,
(	5750	)	,
(	5752	)	,
(	5754	)	,
(	5755	)	,
(	5757	)	,
(	5758	)	,
(	5760	)	,
(	5762	)	,
(	5763	)	,
(	5765	)	,
(	5767	)	,
(	5768	)	,
(	5770	)	,
(	5771	)	,
(	5773	)	,
(	5775	)	,
(	5776	)	,
(	5778	)	,
(	5780	)	,
(	5781	)	,
(	5783	)	,
(	5784	)	,
(	5786	)	,
(	5788	)	,
(	5789	)	,
(	5791	)	,
(	5792	)	,
(	5794	)	,
(	5796	)	,
(	5797	)	,
(	5799	)	,
(	5801	)	,
(	5802	)	,
(	5804	)	,
(	5805	)	,
(	5807	)	,
(	5809	)	,
(	5810	)	,
(	5812	)	,
(	5814	)	,
(	5815	)	,
(	5817	)	,
(	5818	)	,
(	5820	)	,
(	5822	)	,
(	5823	)	,
(	5825	)	,
(	5827	)	,
(	5828	)	,
(	5830	)	,
(	5831	)	,
(	5833	)	,
(	5835	)	,
(	5836	)	,
(	5838	)	,
(	5839	)	,
(	5841	)	,
(	5843	)	,
(	5844	)	,
(	5846	)	,
(	5848	)	,
(	5849	)	,
(	5851	)	,
(	5852	)	,
(	5854	)	,
(	5856	)	,
(	5857	)	,
(	5859	)	,
(	5861	)	,
(	5862	)	,
(	5864	)	,
(	5865	)	,
(	5867	)	,
(	5869	)	,
(	5870	)	,
(	5872	)	,
(	5873	)	,
(	5875	)	,
(	5877	)	,
(	5878	)	,
(	5880	)	,
(	5882	)	,
(	5883	)	,
(	5885	)	,
(	5886	)	,
(	5888	)	,
(	5890	)	,
(	5891	)	,
(	5893	)	,
(	5895	)	,
(	5896	)	,
(	5898	)	,
(	5899	)	,
(	5901	)	,
(	5903	)	,
(	5904	)	,
(	5906	)	,
(	5908	)	,
(	5909	)	,
(	5911	)	,
(	5912	)	,
(	5914	)	,
(	5916	)	,
(	5917	)	,
(	5919	)	,
(	5920	)	,
(	5922	)	,
(	5924	)	,
(	5925	)	,
(	5927	)	,
(	5929	)	,
(	5930	)	,
(	5932	)	,
(	5933	)	,
(	5935	)	,
(	5937	)	,
(	5938	)	,
(	5940	)	,
(	5942	)	,
(	5943	)	,
(	5945	)	,
(	5946	)	,
(	5948	)	,
(	5950	)	,
(	5951	)	,
(	5953	)	,
(	5954	)	,
(	5956	)	,
(	5958	)	,
(	5959	)	,
(	5961	)	,
(	5963	)	,
(	5964	)	,
(	5966	)	,
(	5967	)	,
(	5969	)	,
(	5971	)	,
(	5972	)	,
(	5974	)	,
(	5976	)	,
(	5977	)	,
(	5979	)	,
(	5980	)	,
(	5982	)	,
(	5984	)	,
(	5985	)	,
(	5987	)	,
(	5989	)	,
(	5990	)	,
(	5992	)	,
(	5993	)	,
(	5995	)	,
(	5997	)	,
(	5998	)	,
(	6000	)	,
(	6001	)	,
(	6003	)	,
(	6005	)	,
(	6006	)	,
(	6008	)	,
(	6010	)	,
(	6011	)	,
(	6013	)	,
(	6014	)	,
(	6016	)	,
(	6018	)	,
(	6019	)	,
(	6021	)	,
(	6023	)	,
(	6024	)	,
(	6026	)	,
(	6027	)	,
(	6029	)	,
(	6031	)	,
(	6032	)	,
(	6034	)	,
(	6035	)	,
(	6037	)	,
(	6039	)	,
(	6040	)	,
(	6042	)	,
(	6044	)	,
(	6045	)	,
(	6047	)	,
(	6048	)	,
(	6050	)	,
(	6052	)	,
(	6053	)	,
(	6055	)	,
(	6057	)	,
(	6058	)	,
(	6060	)	,
(	6061	)	,
(	6063	)	,
(	6065	)	,
(	6066	)	,
(	6068	)	,
(	6070	)	,
(	6071	)	,
(	6073	)	,
(	6074	)	,
(	6076	)	,
(	6078	)	,
(	6079	)	,
(	6081	)	,
(	6082	)	,
(	6084	)	,
(	6086	)	,
(	6087	)	,
(	6089	)	,
(	6091	)	,
(	6092	)	,
(	6094	)	,
(	6095	)	,
(	6097	)	,
(	6099	)	,
(	6100	)	,
(	6102	)	,
(	6104	)	,
(	6105	)	,
(	6107	)	,
(	6108	)	,
(	6110	)	,
(	6112	)	,
(	6113	)	,
(	6115	)	,
(	6116	)	,
(	6118	)	,
(	6120	)	,
(	6121	)	,
(	6123	)	,
(	6125	)	,
(	6126	)	,
(	6128	)	,
(	6129	)	,
(	6131	)	,
(	6133	)	,
(	6134	)	,
(	6136	)	,
(	6138	)	,
(	6139	)	,
(	6141	)	,
(	6142	)	,
(	6144	)	,
(	6146	)	,
(	6147	)	,
(	6149	)	,
(	6151	)	,
(	6152	)	,
(	6154	)	,
(	6155	)	,
(	6157	)	,
(	6159	)	,
(	6160	)	,
(	6162	)	,
(	6163	)	,
(	6165	)	,
(	6167	)	,
(	6168	)	,
(	6170	)	,
(	6172	)	,
(	6173	)	,
(	6175	)	,
(	6176	)	,
(	6178	)	,
(	6180	)	,
(	6181	)	,
(	6183	)	,
(	6185	)	,
(	6186	)	,
(	6188	)	,
(	6189	)	,
(	6191	)	,
(	6193	)	,
(	6194	)	,
(	6196	)	,
(	6197	)	,
(	6199	)	,
(	6201	)	,
(	6202	)	,
(	6204	)	,
(	6206	)	,
(	6207	)	,
(	6209	)	,
(	6210	)	,
(	6212	)	,
(	6214	)	,
(	6215	)	,
(	6217	)	,
(	6219	)	,
(	6220	)	,
(	6222	)	,
(	6223	)	,
(	6225	)	,
(	6227	)	,
(	6228	)	,
(	6230	)	,
(	6232	)	,
(	6233	)	,
(	6235	)	,
(	6236	)	,
(	6238	)	,
(	6240	)	,
(	6241	)	,
(	6243	)	,
(	6244	)	,
(	6246	)	,
(	6248	)	,
(	6249	)	,
(	6251	)	,
(	6253	)	,
(	6254	)	,
(	6256	)	,
(	6257	)	,
(	6259	)	,
(	6261	)	,
(	6262	)	,
(	6264	)	,
(	6266	)	,
(	6267	)	,
(	6269	)	,
(	6270	)	,
(	6272	)	,
(	6274	)	,
(	6275	)	,
(	6277	)	,
(	6278	)	,
(	6280	)	,
(	6282	)	,
(	6283	)	,
(	6285	)	,
(	6287	)	,
(	6288	)	,
(	6290	)	,
(	6291	)	,
(	6293	)	,
(	6295	)	,
(	6296	)	,
(	6298	)	,
(	6300	)	,
(	6301	)	,
(	6303	)	,
(	6304	)	,
(	6306	)	,
(	6308	)	,
(	6309	)	,
(	6311	)	,
(	6313	)	,
(	6314	)	,
(	6316	)	,
(	6317	)	,
(	6319	)	,
(	6321	)	,
(	6322	)	,
(	6324	)	,
(	6325	)	,
(	6327	)	,
(	6329	)	,
(	6330	)	,
(	6332	)	,
(	6334	)	,
(	6335	)	,
(	6337	)	,
(	6338	)	,
(	6340	)	,
(	6342	)	,
(	6343	)	,
(	6345	)	,
(	6347	)	,
(	6348	)	,
(	6350	)	,
(	6351	)	,
(	6353	)	,
(	6355	)	,
(	6356	)	,
(	6358	)	,
(	6359	)	,
(	6361	)	,
(	6363	)	,
(	6364	)	,
(	6366	)	,
(	6368	)	,
(	6369	)	,
(	6371	)	,
(	6372	)	,
(	6374	)	,
(	6376	)	,
(	6377	)	,
(	6379	)	,
(	6381	)	,
(	6382	)	,
(	6384	)	,
(	6385	)	,
(	6387	)	,
(	6389	)	,
(	6390	)	,
(	6392	)	,
(	6394	)	,
(	6395	)	,
(	6397	)	,
(	6398	)	,
(	6400	)	,
(	6402	)	,
(	6403	)	,
(	6405	)	,
(	6406	)	,
(	6408	)	,
(	6410	)	,
(	6411	)	,
(	6413	)	,
(	6415	)	,
(	6416	)	,
(	6418	)	,
(	6419	)	,
(	6421	)	,
(	6423	)	,
(	6424	)	,
(	6426	)	,
(	6428	)	,
(	6429	)	,
(	6431	)	,
(	6432	)	,
(	6434	)	,
(	6436	)	,
(	6437	)	,
(	6439	)	,
(	6440	)	,
(	6442	)	,
(	6444	)	,
(	6445	)	,
(	6447	)	,
(	6449	)	,
(	6450	)	,
(	6452	)	,
(	6453	)	,
(	6455	)	,
(	6457	)	,
(	6458	)	,
(	6460	)	,
(	6462	)	,
(	6463	)	,
(	6465	)	,
(	6466	)	,
(	6468	)	,
(	6470	)	,
(	6471	)	,
(	6473	)	,
(	6475	)	,
(	6476	)	,
(	6478	)	,
(	6479	)	,
(	6481	)	,
(	6483	)	,
(	6484	)	,
(	6486	)	,
(	6487	)	,
(	6489	)	,
(	6491	)	,
(	6492	)	,
(	6494	)	,
(	6496	)	,
(	6497	)	,
(	6499	)	,
(	6500	)	,
(	6502	)	,
(	6504	)	,
(	6505	)	,
(	6507	)	,
(	6509	)	,
(	6510	)	,
(	6512	)	,
(	6513	)	,
(	6515	)	,
(	6517	)	,
(	6518	)	,
(	6520	)	,
(	6521	)	,
(	6523	)	,
(	6525	)	,
(	6526	)	,
(	6528	)	,
(	6530	)	,
(	6531	)	,
(	6533	)	,
(	6534	)	,
(	6536	)	,
(	6538	)	,
(	6539	)	,
(	6541	)	,
(	6543	)	,
(	6544	)	,
(	6546	)	,
(	6547	)	,
(	6549	)	,
(	6551	)	,
(	6552	)	,
(	6554	)	,
(	6556	)	,
(	6557	)	,
(	6559	)	,
(	6560	)	,
(	6562	)	,
(	6564	)	,
(	6565	)	,
(	6567	)	,
(	6568	)	,
(	6570	)	,
(	6572	)	,
(	6573	)	,
(	6575	)	,
(	6577	)	,
(	6578	)	,
(	6580	)	,
(	6581	)	,
(	6583	)	,
(	6585	)	,
(	6586	)	,
(	6588	)	,
(	6590	)	,
(	6591	)	,
(	6593	)	,
(	6594	)	,
(	6596	)	,
(	6598	)	,
(	6599	)	,
(	6601	)	,
(	6602	)	,
(	6604	)	,
(	6606	)	,
(	6607	)	,
(	6609	)	,
(	6611	)	,
(	6612	)	,
(	6614	)	,
(	6615	)	,
(	6617	)	,
(	6619	)	,
(	6620	)	,
(	6622	)	,
(	6624	)	,
(	6625	)	,
(	6627	)	,
(	6628	)	,
(	6630	)	,
(	6632	)	,
(	6633	)	,
(	6635	)	,
(	6637	)	,
(	6638	)	,
(	6640	)	,
(	6641	)	,
(	6643	)	,
(	6645	)	,
(	6646	)	,
(	6648	)	,
(	6649	)	,
(	6651	)	,
(	6653	)	,
(	6654	)	,
(	6656	)	,
(	6658	)	,
(	6659	)	,
(	6661	)	,
(	6662	)	,
(	6664	)	,
(	6666	)	,
(	6667	)	,
(	6669	)	,
(	6671	)	,
(	6672	)	,
(	6674	)	,
(	6675	)	,
(	6677	)	,
(	6679	)	,
(	6680	)	,
(	6682	)	,
(	6683	)	,
(	6685	)	,
(	6687	)	,
(	6688	)	,
(	6690	)	,
(	6692	)	,
(	6693	)	,
(	6695	)	,
(	6696	)	,
(	6698	)	,
(	6700	)	,
(	6701	)	,
(	6703	)	,
(	6705	)	,
(	6706	)	,
(	6708	)	,
(	6709	)	,
(	6711	)	,
(	6713	)	,
(	6714	)	,
(	6716	)	,
(	6718	)	,
(	6719	)	,
(	6721	)	,
(	6722	)	,
(	6724	)	,
(	6726	)	,
(	6727	)	,
(	6729	)	,
(	6730	)	,
(	6732	)	,
(	6734	)	,
(	6735	)	,
(	6737	)	,
(	6739	)	,
(	6740	)	,
(	6742	)	,
(	6743	)	,
(	6745	)	,
(	6747	)	,
(	6748	)	,
(	6750	)	,
(	6752	)	,
(	6753	)	,
(	6755	)	,
(	6756	)	,
(	6758	)	,
(	6760	)	,
(	6761	)	,
(	6763	)	,
(	6764	)	,
(	6766	)	,
(	6768	)	,
(	6769	)	,
(	6771	)	,
(	6773	)	,
(	6774	)	,
(	6776	)	,
(	6777	)	,
(	6779	)	,
(	6781	)	,
(	6782	)	,
(	6784	)	,
(	6786	)	,
(	6787	)	,
(	6789	)	,
(	6790	)	,
(	6792	)	,
(	6794	)	,
(	6795	)	,
(	6797	)	,
(	6799	)	,
(	6800	)	,
(	6802	)	,
(	6803	)	,
(	6805	)	,
(	6807	)	,
(	6808	)	,
(	6810	)	,
(	6811	)	,
(	6813	)	,
(	6815	)	,
(	6816	)	,
(	6818	)	,
(	6820	)	,
(	6821	)	,
(	6823	)	,
(	6824	)	,
(	6826	)	,
(	6828	)	,
(	6829	)	,
(	6831	)	,
(	6833	)	,
(	6834	)	,
(	6836	)	,
(	6837	)	,
(	6839	)	,
(	6841	)	,
(	6842	)	,
(	6844	)	,
(	6845	)	,
(	6847	)	,
(	6849	)	,
(	6850	)	,
(	6852	)	,
(	6854	)	,
(	6855	)	,
(	6857	)	,
(	6858	)	,
(	6860	)	,
(	6862	)	,
(	6863	)	,
(	6865	)	,
(	6867	)	,
(	6868	)	,
(	6870	)	,
(	6871	)	,
(	6873	)	,
(	6875	)	,
(	6876	)	,
(	6878	)	,
(	6880	)	,
(	6881	)	,
(	6883	)	,
(	6884	)	,
(	6886	)	,
(	6888	)	,
(	6889	)	,
(	6891	)	,
(	6892	)	,
(	6894	)	,
(	6896	)	,
(	6897	)	,
(	6899	)	,
(	6901	)	,
(	6902	)	,
(	6904	)	,
(	6905	)	,
(	6907	)	,
(	6909	)	,
(	6910	)	,
(	6912	)	,
(	6914	)	,
(	6915	)	,
(	6917	)	,
(	6918	)	,
(	6920	)	,
(	6922	)	,
(	6923	)	,
(	6925	)	,
(	6926	)	,
(	6928	)	,
(	6930	)	,
(	6931	)	,
(	6933	)	,
(	6935	)	,
(	6936	)	,
(	6938	)	,
(	6939	)	,
(	6941	)	,
(	6943	)	,
(	6944	)	,
(	6946	)	,
(	6948	)	,
(	6949	)	,
(	6951	)	,
(	6952	)	,
(	6954	)	,
(	6956	)	,
(	6957	)	,
(	6959	)	,
(	6961	)	,
(	6962	)	,
(	6964	)	,
(	6965	)	,
(	6967	)	,
(	6969	)	,
(	6970	)	,
(	6972	)	,
(	6973	)	,
(	6975	)	,
(	6977	)	,
(	6978	)	,
(	6980	)	,
(	6982	)	,
(	6983	)	,
(	6985	)	,
(	6986	)	,
(	6988	)	,
(	6990	)	,
(	6991	)	,
(	6993	)	,
(	6995	)	,
(	6996	)	,
(	6998	)	,
(	6999	)	,
(	7001	)	,
(	7003	)	,
(	7004	)	,
(	7006	)	,
(	7007	)	,
(	7009	)	,
(	7011	)	,
(	7012	)	,
(	7014	)	,
(	7016	)	,
(	7017	)	,
(	7019	)	,
(	7020	)	,
(	7022	)	,
(	7024	)	,
(	7025	)	,
(	7027	)	,
(	7029	)	,
(	7030	)	,
(	7032	)	,
(	7033	)	,
(	7035	)	,
(	7037	)	,
(	7038	)	,
(	7040	)	,
(	7042	)	,
(	7043	)	,
(	7045	)	,
(	7046	)	,
(	7048	)	,
(	7050	)	,
(	7051	)	,
(	7053	)	,
(	7054	)	,
(	7056	)	,
(	7058	)	,
(	7059	)	,
(	7061	)	,
(	7063	)	,
(	7064	)	,
(	7066	)	,
(	7067	)	,
(	7069	)	,
(	7071	)	,
(	7072	)	,
(	7074	)	,
(	7076	)	,
(	7077	)	,
(	7079	)	,
(	7080	)	,
(	7082	)	,
(	7084	)	,
(	7085	)	,
(	7087	)	,
(	7088	)	,
(	7090	)	,
(	7092	)	,
(	7093	)	,
(	7095	)	,
(	7097	)	,
(	7098	)	,
(	7100	)	,
(	7101	)	,
(	7103	)	,
(	7105	)	,
(	7106	)	,
(	7108	)	,
(	7110	)	,
(	7111	)	,
(	7113	)	,
(	7114	)	,
(	7116	)	,
(	7118	)	,
(	7119	)	,
(	7121	)	,
(	7123	)	,
(	7124	)	,
(	7126	)	,
(	7127	)	,
(	7129	)	,
(	7131	)	,
(	7132	)	,
(	7134	)	,
(	7135	)	,
(	7137	)	,
(	7139	)	,
(	7140	)	,
(	7142	)	,
(	7144	)	,
(	7145	)	,
(	7147	)	,
(	7148	)	,
(	7150	)	,
(	7152	)	,
(	7153	)	,
(	7155	)	,
(	7157	)	,
(	7158	)	,
(	7160	)	,
(	7161	)	,
(	7163	)	,
(	7165	)	,
(	7166	)	,
(	7168	)	,
(	7169	)	,
(	7171	)	,
(	7173	)	,
(	7174	)	,
(	7176	)	,
(	7178	)	,
(	7179	)	,
(	7181	)	,
(	7182	)	,
(	7184	)	,
(	7186	)	,
(	7187	)	,
(	7189	)	,
(	7191	)	,
(	7192	)	,
(	7194	)	,
(	7195	)	,
(	7197	)	,
(	7199	)	,
(	7200	)	,
(	7202	)	,
(	7204	)	,
(	7205	)	,
(	7207	)	,
(	7208	)	,
(	7210	)	,
(	7212	)	,
(	7213	)	,
(	7215	)	,
(	7216	)	,
(	7218	)	,
(	7220	)	,
(	7221	)	,
(	7223	)	,
(	7225	)	,
(	7226	)	,
(	7228	)	,
(	7229	)	,
(	7231	)	,
(	7233	)	,
(	7234	)	,
(	7236	)	,
(	7238	)	,
(	7239	)	,
(	7241	)	,
(	7242	)	,
(	7244	)	,
(	7246	)	,
(	7247	)	,
(	7249	)	,
(	7250	)	,
(	7252	)	,
(	7254	)	,
(	7255	)	,
(	7257	)	,
(	7259	)	,
(	7260	)	,
(	7262	)	,
(	7263	)	,
(	7265	)	,
(	7267	)	,
(	7268	)	,
(	7270	)	,
(	7272	)	,
(	7273	)	,
(	7275	)	,
(	7276	)	,
(	7278	)	,
(	7280	)	,
(	7281	)	,
(	7283	)	,
(	7285	)	,
(	7286	)	,
(	7288	)	,
(	7289	)	,
(	7291	)	,
(	7293	)	,
(	7294	)	,
(	7296	)	,
(	7297	)	,
(	7299	)	,
(	7301	)	,
(	7302	)	,
(	7304	)	,
(	7306	)	,
(	7307	)	,
(	7309	)	,
(	7310	)	,
(	7312	)	,
(	7314	)	,
(	7315	)	,
(	7317	)	,
(	7319	)	,
(	7320	)	,
(	7322	)	,
(	7323	)	,
(	7325	)	,
(	7327	)	,
(	7328	)	,
(	7330	)	,
(	7331	)	,
(	7333	)	,
(	7335	)	,
(	7336	)	,
(	7338	)	,
(	7340	)	,
(	7341	)	,
(	7343	)	,
(	7344	)	,
(	7346	)	,
(	7348	)	,
(	7349	)	,
(	7351	)	,
(	7353	)	,
(	7354	)	,
(	7356	)	,
(	7357	)	,
(	7359	)	,
(	7361	)	,
(	7362	)	,
(	7364	)	,
(	7366	)	,
(	7367	)	,
(	7369	)	,
(	7370	)	,
(	7372	)	,
(	7374	)	,
(	7375	)	,
(	7377	)	,
(	7378	)	,
(	7380	)	,
(	7382	)	,
(	7383	)	,
(	7385	)	,
(	7387	)	,
(	7388	)	,
(	7390	)	,
(	7391	)	,
(	7393	)	,
(	7395	)	,
(	7396	)	,
(	7398	)	,
(	7400	)	,
(	7401	)	,
(	7403	)	,
(	7404	)	,
(	7406	)	,
(	7408	)	,
(	7409	)	,
(	7411	)	,
(	7412	)	,
(	7414	)	,
(	7416	)	,
(	7417	)	,
(	7419	)	,
(	7421	)	,
(	7422	)	,
(	7424	)	,
(	7425	)	,
(	7427	)	,
(	7429	)	,
(	7430	)	,
(	7432	)	,
(	7434	)	,
(	7435	)	,
(	7437	)	,
(	7438	)	,
(	7440	)	,
(	7442	)	,
(	7443	)	,
(	7445	)	,
(	7447	)	,
(	7448	)	,
(	7450	)	,
(	7451	)	,
(	7453	)	,
(	7455	)	,
(	7456	)	,
(	7458	)	,
(	7459	)	,
(	7461	)	,
(	7463	)	,
(	7464	)	,
(	7466	)	,
(	7468	)	,
(	7469	)	,
(	7471	)	,
(	7472	)	,
(	7474	)	,
(	7476	)	,
(	7477	)	,
(	7479	)	,
(	7481	)	,
(	7482	)	,
(	7484	)	,
(	7485	)	,
(	7487	)	,
(	7489	)	,
(	7490	)	,
(	7492	)	,
(	7493	)	,
(	7495	)	,
(	7497	)	,
(	7498	)	,
(	7500	)	,
(	7502	)	,
(	7503	)	,
(	7505	)	,
(	7506	)	,
(	7508	)	,
(	7510	)	,
(	7511	)	,
(	7513	)	,
(	7515	)	,
(	7516	)	,
(	7518	)	,
(	7519	)	,
(	7521	)	,
(	7523	)	,
(	7524	)	,
(	7526	)	,
(	7528	)	,
(	7529	)	,
(	7531	)	,
(	7532	)	,
(	7534	)	,
(	7536	)	,
(	7537	)	,
(	7539	)	,
(	7540	)	,
(	7542	)	,
(	7544	)	,
(	7545	)	,
(	7547	)	,
(	7549	)	,
(	7550	)	,
(	7552	)	,
(	7553	)	,
(	7555	)	,
(	7557	)	,
(	7558	)	,
(	7560	)	,
(	7562	)	,
(	7563	)	,
(	7565	)	,
(	7566	)	,
(	7568	)	,
(	7570	)	,
(	7571	)	,
(	7573	)	,
(	7574	)	,
(	7576	)	,
(	7578	)	,
(	7579	)	,
(	7581	)	,
(	7583	)	,
(	7584	)	,
(	7586	)	,
(	7587	)	,
(	7589	)	,
(	7591	)	,
(	7592	)	,
(	7594	)	,
(	7596	)	,
(	7597	)	,
(	7599	)	,
(	7600	)	,
(	7602	)	,
(	7604	)	,
(	7605	)	,
(	7607	)	,
(	7609	)	,
(	7610	)	,
(	7612	)	,
(	7613	)	,
(	7615	)	,
(	7617	)	,
(	7618	)	,
(	7620	)	,
(	7621	)	,
(	7623	)	,
(	7625	)	,
(	7626	)	,
(	7628	)	,
(	7630	)	,
(	7631	)	,
(	7633	)	,
(	7634	)	,
(	7636	)	,
(	7638	)	,
(	7639	)	,
(	7641	)	,
(	7643	)	,
(	7644	)	,
(	7646	)	,
(	7647	)	,
(	7649	)	,
(	7651	)	,
(	7652	)	,
(	7654	)	,
(	7655	)	,
(	7657	)	,
(	7659	)	,
(	7660	)	,
(	7662	)	,
(	7664	)	,
(	7665	)	,
(	7667	)	,
(	7668	)	,
(	7670	)	,
(	7672	)	,
(	7673	)	,
(	7675	)	,
(	7677	)	,
(	7678	)	,
(	7680	)	,
(	7681	)	,
(	7683	)	,
(	7685	)	,
(	7686	)	,
(	7688	)	,
(	7690	)	,
(	7691	)	,
(	7693	)	,
(	7694	)	,
(	7696	)	,
(	7698	)	,
(	7699	)	,
(	7701	)	,
(	7702	)	,
(	7704	)	,
(	7706	)	,
(	7707	)	,
(	7709	)	,
(	7711	)	,
(	7712	)	,
(	7714	)	,
(	7715	)	,
(	7717	)	,
(	7719	)	,
(	7720	)	,
(	7722	)	,
(	7724	)	,
(	7725	)	,
(	7727	)	,
(	7728	)	,
(	7730	)	,
(	7732	)	,
(	7733	)	,
(	7735	)	,
(	7736	)	,
(	7738	)	,
(	7740	)	,
(	7741	)	,
(	7743	)	,
(	7745	)	,
(	7746	)	,
(	7748	)	,
(	7749	)	,
(	7751	)	,
(	7753	)	,
(	7754	)	,
(	7756	)	,
(	7758	)	,
(	7759	)	,
(	7761	)	,
(	7762	)	,
(	7764	)	,
(	7766	)	,
(	7767	)	,
(	7769	)	,
(	7771	)	,
(	7772	)	,
(	7774	)	,
(	7775	)	,
(	7777	)	,
(	7779	)	,
(	7780	)	,
(	7782	)	,
(	7783	)	,
(	7785	)	,
(	7787	)	,
(	7788	)	,
(	7790	)	,
(	7792	)	,
(	7793	)	,
(	7795	)	,
(	7796	)	,
(	7798	)	,
(	7800	)	,
(	7801	)	,
(	7803	)	,
(	7805	)	,
(	7806	)	,
(	7808	)	,
(	7809	)	,
(	7811	)	,
(	7813	)	,
(	7814	)	,
(	7816	)	,
(	7817	)	,
(	7819	)	,
(	7821	)	,
(	7822	)	,
(	7824	)	,
(	7826	)	,
(	7827	)	,
(	7829	)	,
(	7830	)	,
(	7832	)	,
(	7834	)	,
(	7835	)	,
(	7837	)	,
(	7839	)	,
(	7840	)	,
(	7842	)	,
(	7843	)	,
(	7845	)	,
(	7847	)	,
(	7848	)	,
(	7850	)	,
(	7852	)	,
(	7853	)	,
(	7855	)	,
(	7856	)	,
(	7858	)	,
(	7860	)	,
(	7861	)	,
(	7863	)	,
(	7864	)	,
(	7866	)	,
(	7868	)	,
(	7869	)	,
(	7871	)	,
(	7873	)	,
(	7874	)	,
(	7876	)	,
(	7877	)	,
(	7879	)	,
(	7881	)	,
(	7882	)	,
(	7884	)	,
(	7886	)	,
(	7887	)	,
(	7889	)	,
(	7890	)	,
(	7892	)	,
(	7894	)	,
(	7895	)	,
(	7897	)	,
(	7898	)	,
(	7900	)	,
(	7902	)	,
(	7903	)	,
(	7905	)	,
(	7907	)	,
(	7908	)	,
(	7910	)	,
(	7911	)	,
(	7913	)	,
(	7915	)	,
(	7916	)	,
(	7918	)	,
(	7920	)	,
(	7921	)	,
(	7923	)	,
(	7924	)	,
(	7926	)	,
(	7928	)	,
(	7929	)	,
(	7931	)	,
(	7933	)	,
(	7934	)	,
(	7936	)	,
(	7937	)	,
(	7939	)	,
(	7941	)	,
(	7942	)	,
(	7944	)	,
(	7945	)	,
(	7947	)	,
(	7949	)	,
(	7950	)	,
(	7952	)	,
(	7954	)	,
(	7955	)	,
(	7957	)	,
(	7958	)	,
(	7960	)	,
(	7962	)	,
(	7963	)	,
(	7965	)	,
(	7967	)	,
(	7968	)	,
(	7970	)	,
(	7971	)	,
(	7973	)	,
(	7975	)	,
(	7976	)	,
(	7978	)	,
(	7979	)	,
(	7981	)	,
(	7983	)	,
(	7984	)	,
(	7986	)	,
(	7988	)	,
(	7989	)	,
(	7991	)	,
(	7992	)	,
(	7994	)	,
(	7996	)	,
(	7997	)	,
(	7999	)	,
(	8001	)	,
(	8002	)	,
(	8004	)	,
(	8005	)	,
(	8007	)	,
(	8009	)	,
(	8010	)	,
(	8012	)	,
(	8014	)	,
(	8015	)	,
(	8017	)	,
(	8018	)	,
(	8020	)	,
(	8022	)	,
(	8023	)	,
(	8025	)	,
(	8026	)	,
(	8028	)	,
(	8030	)	,
(	8031	)	,
(	8033	)	,
(	8035	)	,
(	8036	)	,
(	8038	)	,
(	8039	)	,
(	8041	)	,
(	8043	)	,
(	8044	)	,
(	8046	)	,
(	8048	)	,
(	8049	)	,
(	8051	)	,
(	8052	)	,
(	8054	)	,
(	8056	)	,
(	8057	)	,
(	8059	)	,
(	8060	)	,
(	8062	)	,
(	8064	)	,
(	8065	)	,
(	8067	)	,
(	8069	)	,
(	8070	)	,
(	8072	)	,
(	8073	)	,
(	8075	)	,
(	8077	)	,
(	8078	)	,
(	8080	)	,
(	8082	)	,
(	8083	)	,
(	8085	)	,
(	8086	)	,
(	8088	)	,
(	8090	)	,
(	8091	)	,
(	8093	)	,
(	8095	)	,
(	8096	)	,
(	8098	)	,
(	8099	)	,
(	8101	)	,
(	8103	)	,
(	8104	)	,
(	8106	)	,
(	8107	)	,
(	8109	)	,
(	8111	)	,
(	8112	)	,
(	8114	)	,
(	8116	)	,
(	8117	)	,
(	8119	)	,
(	8120	)	,
(	8122	)	,
(	8124	)	,
(	8125	)	,
(	8127	)	,
(	8129	)	,
(	8130	)	,
(	8132	)	,
(	8133	)	,
(	8135	)	,
(	8137	)	,
(	8138	)	,
(	8140	)	,
(	8141	)	,
(	8143	)	,
(	8145	)	,
(	8146	)	,
(	8148	)	,
(	8150	)	,
(	8151	)	,
(	8153	)	,
(	8154	)	,
(	8156	)	,
(	8158	)	,
(	8159	)	,
(	8161	)	,
(	8163	)	,
(	8164	)	,
(	8166	)	,
(	8167	)	,
(	8169	)	,
(	8171	)	,
(	8172	)	,
(	8174	)	,
(	8176	)	,
(	8177	)	,
(	8179	)	,
(	8180	)	,
(	8182	)	,
(	8184	)	,
(	8185	)	,
(	8187	)	,
(	8188	)	,
(	8190	)	,
(	8192	)	,
(	8193	)	,
(	8195	)	,
(	8197	)	,
(	8198	)	,
(	8200	)	,
(	8201	)	,
(	8203	)	,
(	8205	)	,
(	8206	)	,
(	8208	)	,
(	8210	)	,
(	8211	)	,
(	8213	)	,
(	8214	)	,
(	8216	)	,
(	8218	)	,
(	8219	)	,
(	8221	)	,
(	8222	)	,
(	8224	)	,
(	8226	)	,
(	8227	)	,
(	8229	)	,
(	8231	)	,
(	8232	)	,
(	8234	)	,
(	8235	)	,
(	8237	)	,
(	8239	)	,
(	8240	)	,
(	8242	)	,
(	8244	)	,
(	8245	)	,
(	8247	)	,
(	8248	)	,
(	8250	)	,
(	8252	)	,
(	8253	)	,
(	8255	)	,
(	8257	)	,
(	8258	)	,
(	8260	)	,
(	8261	)	,
(	8263	)	,
(	8265	)	,
(	8266	)	,
(	8268	)	,
(	8269	)	,
(	8271	)	,
(	8273	)	,
(	8274	)	,
(	8276	)	,
(	8278	)	,
(	8279	)	,
(	8281	)	,
(	8282	)	,
(	8284	)	,
(	8286	)	,
(	8287	)	,
(	8289	)	,
(	8291	)	,
(	8292	)	,
(	8294	)	,
(	8295	)	,
(	8297	)	,
(	8299	)	,
(	8300	)	,
(	8302	)	,
(	8303	)	,
(	8305	)	,
(	8307	)	,
(	8308	)	,
(	8310	)	,
(	8312	)	,
(	8313	)	,
(	8315	)	,
(	8316	)	,
(	8318	)	,
(	8320	)	,
(	8321	)	,
(	8323	)	,
(	8325	)	,
(	8326	)	,
(	8328	)	,
(	8329	)	,
(	8331	)	,
(	8333	)	,
(	8334	)	,
(	8336	)	,
(	8338	)	,
(	8339	)	,
(	8341	)	,
(	8342	)	,
(	8344	)	,
(	8346	)	,
(	8347	)	,
(	8349	)	,
(	8350	)	,
(	8352	)	,
(	8354	)	,
(	8355	)	,
(	8357	)	,
(	8359	)	,
(	8360	)	,
(	8362	)	,
(	8363	)	,
(	8365	)	,
(	8367	)	,
(	8368	)	,
(	8370	)	,
(	8372	)	,
(	8373	)	,
(	8375	)	,
(	8376	)	,
(	8378	)	,
(	8380	)	,
(	8381	)	,
(	8383	)	,
(	8384	)	,
(	8386	)	,
(	8388	)	,
(	8389	)	,
(	8391	)	,
(	8393	)	,
(	8394	)	,
(	8396	)	,
(	8397	)	,
(	8399	)	,
(	8401	)	,
(	8402	)	,
(	8404	)	,
(	8406	)	,
(	8407	)	,
(	8409	)	,
(	8410	)	,
(	8412	)	,
(	8414	)	,
(	8415	)	,
(	8417	)	,
(	8419	)	,
(	8420	)	,
(	8422	)	,
(	8423	)	,
(	8425	)	,
(	8427	)	,
(	8428	)	,
(	8430	)	,
(	8431	)	,
(	8433	)	,
(	8435	)	,
(	8436	)	,
(	8438	)	,
(	8440	)	,
(	8441	)	,
(	8443	)	,
(	8444	)	,
(	8446	)	,
(	8448	)	,
(	8449	)	,
(	8451	)	,
(	8453	)	,
(	8454	)	,
(	8456	)	,
(	8457	)	,
(	8459	)	,
(	8461	)	,
(	8462	)	,
(	8464	)	,
(	8465	)	,
(	8467	)	,
(	8469	)	,
(	8470	)	,
(	8472	)	,
(	8474	)	,
(	8475	)	,
(	8477	)	,
(	8478	)	,
(	8480	)	,
(	8482	)	,
(	8483	)	,
(	8485	)	,
(	8487	)	,
(	8488	)	,
(	8490	)	,
(	8491	)	,
(	8493	)	,
(	8495	)	,
(	8496	)	,
(	8498	)	,
(	8500	)	,
(	8501	)	,
(	8503	)	,
(	8504	)	,
(	8506	)	,
(	8508	)	,
(	8509	)	,
(	8511	)	,
(	8512	)	,
(	8514	)	,
(	8516	)	,
(	8517	)	,
(	8519	)	,
(	8521	)	,
(	8522	)	,
(	8524	)	,
(	8525	)	,
(	8527	)	,
(	8529	)	,
(	8530	)	,
(	8532	)	,
(	8534	)	,
(	8535	)	,
(	8537	)	,
(	8538	)	,
(	8540	)	,
(	8542	)	,
(	8543	)	,
(	8545	)	,
(	8546	)	,
(	8548	)	,
(	8550	)	,
(	8551	)	,
(	8553	)	,
(	8555	)	,
(	8556	)	,
(	8558	)	,
(	8559	)	,
(	8561	)	,
(	8563	)	,
(	8564	)	,
(	8566	)	,
(	8568	)	,
(	8569	)	,
(	8571	)	,
(	8572	)	,
(	8574	)	,
(	8576	)	,
(	8577	)	,
(	8579	)	,
(	8581	)	,
(	8582	)	,
(	8584	)	,
(	8585	)	,
(	8587	)	,
(	8589	)	,
(	8590	)	,
(	8592	)	,
(	8593	)	,
(	8595	)	,
(	8597	)	,
(	8598	)	,
(	8600	)	,
(	8602	)	,
(	8603	)	,
(	8605	)	,
(	8606	)	,
(	8608	)	,
(	8610	)	,
(	8611	)	,
(	8613	)	,
(	8615	)	,
(	8616	)	,
(	8618	)	,
(	8619	)	,
(	8621	)	,
(	8623	)	,
(	8624	)	,
(	8626	)	,
(	8627	)	,
(	8629	)	,
(	8631	)	,
(	8632	)	,
(	8634	)	,
(	8636	)	,
(	8637	)	,
(	8639	)	,
(	8640	)	,
(	8642	)	,
(	8644	)	,
(	8645	)	,
(	8647	)	,
(	8649	)	,
(	8650	)	,
(	8652	)	,
(	8653	)	,
(	8655	)	,
(	8657	)	,
(	8658	)	,
(	8660	)	,
(	8662	)	,
(	8663	)	,
(	8665	)	,
(	8666	)	,
(	8668	)	,
(	8670	)	,
(	8671	)	,
(	8673	)	,
(	8674	)	,
(	8676	)	,
(	8678	)	,
(	8679	)	,
(	8681	)	,
(	8683	)	,
(	8684	)	,
(	8686	)	,
(	8687	)	,
(	8689	)	,
(	8691	)	,
(	8692	)	,
(	8694	)	,
(	8696	)	,
(	8697	)	,
(	8699	)	,
(	8700	)	,
(	8702	)	,
(	8704	)	,
(	8705	)	,
(	8707	)	,
(	8708	)	,
(	8710	)	,
(	8712	)	,
(	8713	)	,
(	8715	)	,
(	8717	)	,
(	8718	)	,
(	8720	)	,
(	8721	)	,
(	8723	)	,
(	8725	)	,
(	8726	)	,
(	8728	)	,
(	8730	)	,
(	8731	)	,
(	8733	)	,
(	8734	)	,
(	8736	)	,
(	8738	)	,
(	8739	)	,
(	8741	)	,
(	8743	)	,
(	8744	)	,
(	8746	)	,
(	8747	)	,
(	8749	)	,
(	8751	)	,
(	8752	)	,
(	8754	)	,
(	8755	)	,
(	8757	)	,
(	8759	)	,
(	8760	)	,
(	8762	)	,
(	8764	)	,
(	8765	)	,
(	8767	)	,
(	8768	)	,
(	8770	)	,
(	8772	)	,
(	8773	)	,
(	8775	)	,
(	8777	)	,
(	8778	)	,
(	8780	)	,
(	8781	)	,
(	8783	)	,
(	8785	)	,
(	8786	)	,
(	8788	)	,
(	8789	)	,
(	8791	)	,
(	8793	)	,
(	8794	)	,
(	8796	)	,
(	8798	)	,
(	8799	)	,
(	8801	)	,
(	8802	)	,
(	8804	)	,
(	8806	)	,
(	8807	)	,
(	8809	)	,
(	8811	)	,
(	8812	)	,
(	8814	)	,
(	8815	)	,
(	8817	)	,
(	8819	)	,
(	8820	)	,
(	8822	)	,
(	8824	)	,
(	8825	)	,
(	8827	)	,
(	8828	)	,
(	8830	)	,
(	8832	)	,
(	8833	)	,
(	8835	)	,
(	8836	)	,
(	8838	)	,
(	8840	)	,
(	8841	)	,
(	8843	)	,
(	8845	)	,
(	8846	)	,
(	8848	)	,
(	8849	)	,
(	8851	)	,
(	8853	)	,
(	8854	)	,
(	8856	)	,
(	8858	)	,
(	8859	)	,
(	8861	)	,
(	8862	)	,
(	8864	)	,
(	8866	)	,
(	8867	)	,
(	8869	)	,
(	8870	)	,
(	8872	)	,
(	8874	)	,
(	8875	)	,
(	8877	)	,
(	8879	)	,
(	8880	)	,
(	8882	)	,
(	8883	)	,
(	8885	)	,
(	8887	)	,
(	8888	)	,
(	8890	)	,
(	8892	)	,
(	8893	)	,
(	8895	)	,
(	8896	)	,
(	8898	)	,
(	8900	)	,
(	8901	)	,
(	8903	)	,
(	8905	)	,
(	8906	)	,
(	8908	)	,
(	8909	)	,
(	8911	)	,
(	8913	)	,
(	8914	)	,
(	8916	)	,
(	8917	)	,
(	8919	)	,
(	8921	)	,
(	8922	)	,
(	8924	)	,
(	8926	)	,
(	8927	)	,
(	8929	)	,
(	8930	)	,
(	8932	)	,
(	8934	)	,
(	8935	)	,
(	8937	)	,
(	8939	)	,
(	8940	)	,
(	8942	)	,
(	8943	)	,
(	8945	)	,
(	8947	)	,
(	8948	)	,
(	8950	)	,
(	8951	)	,
(	8953	)	,
(	8955	)	,
(	8956	)	,
(	8958	)	,
(	8960	)	,
(	8961	)	,
(	8963	)	,
(	8964	)	,
(	8966	)	,
(	8968	)	,
(	8969	)	,
(	8971	)	,
(	8973	)	,
(	8974	)	,
(	8976	)	,
(	8977	)	,
(	8979	)	,
(	8981	)	,
(	8982	)	,
(	8984	)	,
(	8986	)	,
(	8987	)	,
(	8989	)	,
(	8990	)	,
(	8992	)	,
(	8994	)	,
(	8995	)	,
(	8997	)	,
(	8998	)	,
(	9000	)	,
(	9002	)	,
(	9003	)	,
(	9005	)	,
(	9007	)	,
(	9008	)	,
(	9010	)	,
(	9011	)	,
(	9013	)	,
(	9015	)	,
(	9016	)	,
(	9018	)	,
(	9020	)	,
(	9021	)	,
(	9023	)	,
(	9024	)	,
(	9026	)	,
(	9028	)	,
(	9029	)	,
(	9031	)	,
(	9032	)	,
(	9034	)	,
(	9036	)	,
(	9037	)	,
(	9039	)	,
(	9041	)	,
(	9042	)	,
(	9044	)	,
(	9045	)	,
(	9047	)	,
(	9049	)	,
(	9050	)	,
(	9052	)	,
(	9054	)	,
(	9055	)	,
(	9057	)	,
(	9058	)	,
(	9060	)	,
(	9062	)	,
(	9063	)	,
(	9065	)	,
(	9067	)	,
(	9068	)	,
(	9070	)	,
(	9071	)	,
(	9073	)	,
(	9075	)	,
(	9076	)	,
(	9078	)	,
(	9079	)	,
(	9081	)	,
(	9083	)	,
(	9084	)	,
(	9086	)	,
(	9088	)	,
(	9089	)	,
(	9091	)	,
(	9092	)	,
(	9094	)	,
(	9096	)	,
(	9097	)	,
(	9099	)	,
(	9101	)	,
(	9102	)	,
(	9104	)	,
(	9105	)	,
(	9107	)	,
(	9109	)	,
(	9110	)	,
(	9112	)	,
(	9113	)	,
(	9115	)	,
(	9117	)	,
(	9118	)	,
(	9120	)	,
(	9122	)	,
(	9123	)	,
(	9125	)	,
(	9126	)	,
(	9128	)	,
(	9130	)	,
(	9131	)	,
(	9133	)	,
(	9135	)	,
(	9136	)	,
(	9138	)	,
(	9139	)	,
(	9141	)	,
(	9143	)	,
(	9144	)	,
(	9146	)	,
(	9148	)	,
(	9149	)	,
(	9151	)	,
(	9152	)	,
(	9154	)	,
(	9156	)	,
(	9157	)	,
(	9159	)	,
(	9160	)	,
(	9162	)	,
(	9164	)	,
(	9165	)	,
(	9167	)	,
(	9169	)	,
(	9170	)	,
(	9172	)	,
(	9173	)	,
(	9175	)	,
(	9177	)	,
(	9178	)	,
(	9180	)	,
(	9182	)	,
(	9183	)	,
(	9185	)	,
(	9186	)	,
(	9188	)	,
(	9190	)	,
(	9191	)	,
(	9193	)	,
(	9194	)	,
(	9196	)	,
(	9198	)	,
(	9199	)	,
(	9201	)	,
(	9203	)	,
(	9204	)	,
(	9206	)	,
(	9207	)	,
(	9209	)	,
(	9211	)	,
(	9212	)	,
(	9214	)	,
(	9216	)	,
(	9217	)	,
(	9219	)	,
(	9220	)	,
(	9222	)	,
(	9224	)	,
(	9225	)	,
(	9227	)	,
(	9229	)	,
(	9230	)	,
(	9232	)	,
(	9233	)	,
(	9235	)	,
(	9237	)	,
(	9238	)	,
(	9240	)	,
(	9241	)	,
(	9243	)	,
(	9245	)	,
(	9246	)	,
(	9248	)	,
(	9250	)	,
(	9251	)	,
(	9253	)	,
(	9254	)	,
(	9256	)	,
(	9258	)	,
(	9259	)	,
(	9261	)	,
(	9263	)	,
(	9264	)	,
(	9266	)	,
(	9267	)	,
(	9269	)	,
(	9271	)	,
(	9272	)	,
(	9274	)	,
(	9275	)	,
(	9277	)	,
(	9279	)	,
(	9280	)	,
(	9282	)	,
(	9284	)	,
(	9285	)	,
(	9287	)	,
(	9288	)	,
(	9290	)	,
(	9292	)	,
(	9293	)	,
(	9295	)	,
(	9297	)	,
(	9298	)	,
(	9300	)	,
(	9301	)	,
(	9303	)	,
(	9305	)	,
(	9306	)	,
(	9308	)	,
(	9310	)	,
(	9311	)	,
(	9313	)	,
(	9314	)	,
(	9316	)	,
(	9318	)	,
(	9319	)	,
(	9321	)	,
(	9322	)	,
(	9324	)	,
(	9326	)	,
(	9327	)	,
(	9329	)	,
(	9331	)	,
(	9332	)	,
(	9334	)	,
(	9335	)	,
(	9337	)	,
(	9339	)	,
(	9340	)	,
(	9342	)	,
(	9344	)	,
(	9345	)	,
(	9347	)	,
(	9348	)	,
(	9350	)	,
(	9352	)	,
(	9353	)	,
(	9355	)	,
(	9356	)	,
(	9358	)	,
(	9360	)	,
(	9361	)	,
(	9363	)	,
(	9365	)	,
(	9366	)	,
(	9368	)	,
(	9369	)	,
(	9371	)	,
(	9373	)	,
(	9374	)	,
(	9376	)	,
(	9378	)	,
(	9379	)	,
(	9381	)	,
(	9382	)	,
(	9384	)	,
(	9386	)	,
(	9387	)	,
(	9389	)	,
(	9391	)	,
(	9392	)	,
(	9394	)	,
(	9395	)	,
(	9397	)	,
(	9399	)	,
(	9400	)	,
(	9402	)	,
(	9403	)	,
(	9405	)	,
(	9407	)	,
(	9408	)	,
(	9410	)	,
(	9412	)	,
(	9413	)	,
(	9415	)	,
(	9416	)	,
(	9418	)	,
(	9420	)	,
(	9421	)	,
(	9423	)	,
(	9425	)	,
(	9426	)	,
(	9428	)	,
(	9429	)	,
(	9431	)	,
(	9433	)	,
(	9434	)	,
(	9436	)	,
(	9437	)	,
(	9439	)	,
(	9441	)	,
(	9442	)	,
(	9444	)	,
(	9446	)	,
(	9447	)	,
(	9449	)	,
(	9450	)	,
(	9452	)	,
(	9454	)	,
(	9455	)	,
(	9457	)	,
(	9459	)	,
(	9460	)	,
(	9462	)	,
(	9463	)	,
(	9465	)	,
(	9467	)	,
(	9468	)	,
(	9470	)	,
(	9472	)	,
(	9473	)	,
(	9475	)	,
(	9476	)	,
(	9478	)	,
(	9480	)	,
(	9481	)	,
(	9483	)	,
(	9484	)	,
(	9486	)	,
(	9488	)	,
(	9489	)	,
(	9491	)	,
(	9493	)	,
(	9494	)	,
(	9496	)	,
(	9497	)	,
(	9499	)	,
(	9501	)	,
(	9502	)	,
(	9504	)	,
(	9506	)	,
(	9507	)	,
(	9509	)	,
(	9510	)	,
(	9512	)	,
(	9514	)	,
(	9515	)	,
(	9517	)	,
(	9518	)	,
(	9520	)	,
(	9522	)	,
(	9523	)	,
(	9525	)	,
(	9527	)	,
(	9528	)	,
(	9530	)	,
(	9531	)	,
(	9533	)	,
(	9535	)	,
(	9536	)	,
(	9538	)	,
(	9540	)	,
(	9541	)	,
(	9543	)	,
(	9544	)	,
(	9546	)	,
(	9548	)	,
(	9549	)	,
(	9551	)	,
(	9553	)	,
(	9554	)	,
(	9556	)	,
(	9557	)	,
(	9559	)	,
(	9561	)	,
(	9562	)	,
(	9564	)	,
(	9565	)	,
(	9567	)	,
(	9569	)	,
(	9570	)	,
(	9572	)	,
(	9574	)	,
(	9575	)	,
(	9577	)	,
(	9578	)	,
(	9580	)	,
(	9582	)	,
(	9583	)	,
(	9585	)	,
(	9587	)	,
(	9588	)	,
(	9590	)	,
(	9591	)	,
(	9593	)	,
(	9595	)	,
(	9596	)	,
(	9598	)	,
(	9599	)	,
(	9601	)	,
(	9603	)	,
(	9604	)	,
(	9606	)	,
(	9608	)	,
(	9609	)	,
(	9611	)	,
(	9612	)	,
(	9614	)	,
(	9616	)	,
(	9617	)	,
(	9619	)	,
(	9621	)	,
(	9622	)	,
(	9624	)	,
(	9625	)	,
(	9627	)	,
(	9629	)	,
(	9630	)	,
(	9632	)	,
(	9634	)	,
(	9635	)	,
(	9637	)	,
(	9638	)	,
(	9640	)	,
(	9642	)	,
(	9643	)	,
(	9645	)	,
(	9646	)	,
(	9648	)	,
(	9650	)	,
(	9651	)	,
(	9653	)	,
(	9655	)	,
(	9656	)	,
(	9658	)	,
(	9659	)	,
(	9661	)	,
(	9663	)	,
(	9664	)	,
(	9666	)	,
(	9668	)	,
(	9669	)	,
(	9671	)	,
(	9672	)	,
(	9674	)	,
(	9676	)	,
(	9677	)	,
(	9679	)	,
(	9680	)	,
(	9682	)	,
(	9684	)	,
(	9685	)	,
(	9687	)	,
(	9689	)	,
(	9690	)	,
(	9692	)	,
(	9693	)	,
(	9695	)	,
(	9697	)	,
(	9698	)	,
(	9700	)	,
(	9702	)	,
(	9703	)	,
(	9705	)	,
(	9706	)	,
(	9708	)	,
(	9710	)	,
(	9711	)	,
(	9713	)	,
(	9715	)	,
(	9716	)	,
(	9718	)	,
(	9719	)	,
(	9721	)	,
(	9723	)	,
(	9724	)	,
(	9726	)	,
(	9727	)	,
(	9729	)	,
(	9731	)	,
(	9732	)	,
(	9734	)	,
(	9736	)	,
(	9737	)	,
(	9739	)	,
(	9740	)	,
(	9742	)	,
(	9744	)	,
(	9745	)	,
(	9747	)	,
(	9749	)	,
(	9750	)	,
(	9752	)	,
(	9753	)	,
(	9755	)	,
(	9757	)	,
(	9758	)	,
(	9760	)	,
(	9761	)	,
(	9763	)	,
(	9765	)	,
(	9766	)	,
(	9768	)	,
(	9770	)	,
(	9771	)	,
(	9773	)	,
(	9774	)	,
(	9776	)	,
(	9778	)	,
(	9779	)	,
(	9781	)	,
(	9783	)	,
(	9784	)	,
(	9786	)	,
(	9787	)	,
(	9789	)	,
(	9791	)	,
(	9792	)	,
(	9794	)	,
(	9796	)	,
(	9797	)	,
(	9799	)	,
(	9800	)	,
(	9802	)	,
(	9804	)	,
(	9805	)	,
(	9807	)	,
(	9808	)	,
(	9810	)	,
(	9812	)	,
(	9813	)	,
(	9815	)	,
(	9817	)	,
(	9818	)	,
(	9820	)	,
(	9821	)	,
(	9823	)	,
(	9825	)	,
(	9826	)	,
(	9828	)	,
(	9830	)	,
(	9831	)	,
(	9833	)	,
(	9834	)	,
(	9836	)	,
(	9838	)	,
(	9839	)	,
(	9841	)	,
(	9842	)	,
(	9844	)	,
(	9846	)	,
(	9847	)	,
(	9849	)	,
(	9851	)	,
(	9852	)	,
(	9854	)	,
(	9855	)	,
(	9857	)	,
(	9859	)	,
(	9860	)	,
(	9862	)	,
(	9864	)	,
(	9865	)	,
(	9867	)	,
(	9868	)	,
(	9870	)	,
(	9872	)	,
(	9873	)	,
(	9875	)	,
(	9877	)	,
(	9878	)	,
(	9880	)	,
(	9881	)	,
(	9883	)	,
(	9885	)	,
(	9886	)	,
(	9888	)	,
(	9889	)	,
(	9891	)	,
(	9893	)	,
(	9894	)	,
(	9896	)	,
(	9898	)	,
(	9899	)	,
(	9901	)	,
(	9902	)	,
(	9904	)	,
(	9906	)	,
(	9907	)	,
(	9909	)	,
(	9911	)	,
(	9912	)	,
(	9914	)	,
(	9915	)	,
(	9917	)	,
(	9919	)	,
(	9920	)	,
(	9922	)	,
(	9923	)	,
(	9925	)	,
(	9927	)	,
(	9928	)	,
(	9930	)	,
(	9932	)	,
(	9933	)	,
(	9935	)	,
(	9936	)	,
(	9938	)	,
(	9940	)	,
(	9941	)	,
(	9943	)	,
(	9945	)	,
(	9946	)	,
(	9948	)	,
(	9949	)	,
(	9951	)	,
(	9953	)	,
(	9954	)	,
(	9956	)	,
(	9958	)	,
(	9959	)	,
(	9961	)	,
(	9962	)	,
(	9964	)	,
(	9966	)	,
(	9967	)	
						-- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
    	
   frequency <= v2f_LUT(to_integer(unsigned(voltage)));

end behavior;
