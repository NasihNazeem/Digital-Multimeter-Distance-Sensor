LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2frequency IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      frequency      :  OUT   natural
		);		
END voltage2frequency;

ARCHITECTURE behavior OF voltage2frequency IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are maximum counters that will be input
-- into PWM_DAC. The equation used to map a distance to a frequency
-- can be found in an excel (voltage2frequency.xls) file.

type array_1d is array (0 to 4095) of integer;
constant v2f_LUT : array_1d := (

(	10000	)	,
(	9998	)	,
(	9997	)	,
(	9995	)	,
(	9994	)	,
(	9992	)	,
(	9990	)	,
(	9989	)	,
(	9987	)	,
(	9985	)	,
(	9984	)	,
(	9982	)	,
(	9981	)	,
(	9979	)	,
(	9977	)	,
(	9976	)	,
(	9974	)	,
(	9972	)	,
(	9971	)	,
(	9969	)	,
(	9968	)	,
(	9966	)	,
(	9964	)	,
(	9963	)	,
(	9961	)	,
(	9959	)	,
(	9958	)	,
(	9956	)	,
(	9955	)	,
(	9953	)	,
(	9951	)	,
(	9950	)	,
(	9948	)	,
(	9947	)	,
(	9945	)	,
(	9943	)	,
(	9942	)	,
(	9940	)	,
(	9938	)	,
(	9937	)	,
(	9935	)	,
(	9934	)	,
(	9932	)	,
(	9930	)	,
(	9929	)	,
(	9927	)	,
(	9925	)	,
(	9924	)	,
(	9922	)	,
(	9921	)	,
(	9919	)	,
(	9917	)	,
(	9916	)	,
(	9914	)	,
(	9913	)	,
(	9911	)	,
(	9909	)	,
(	9908	)	,
(	9906	)	,
(	9904	)	,
(	9903	)	,
(	9901	)	,
(	9900	)	,
(	9898	)	,
(	9896	)	,
(	9895	)	,
(	9893	)	,
(	9891	)	,
(	9890	)	,
(	9888	)	,
(	9887	)	,
(	9885	)	,
(	9883	)	,
(	9882	)	,
(	9880	)	,
(	9878	)	,
(	9877	)	,
(	9875	)	,
(	9874	)	,
(	9872	)	,
(	9870	)	,
(	9869	)	,
(	9867	)	,
(	9866	)	,
(	9864	)	,
(	9862	)	,
(	9861	)	,
(	9859	)	,
(	9857	)	,
(	9856	)	,
(	9854	)	,
(	9853	)	,
(	9851	)	,
(	9849	)	,
(	9848	)	,
(	9846	)	,
(	9844	)	,
(	9843	)	,
(	9841	)	,
(	9840	)	,
(	9838	)	,
(	9836	)	,
(	9835	)	,
(	9833	)	,
(	9832	)	,
(	9830	)	,
(	9828	)	,
(	9827	)	,
(	9825	)	,
(	9823	)	,
(	9822	)	,
(	9820	)	,
(	9819	)	,
(	9817	)	,
(	9815	)	,
(	9814	)	,
(	9812	)	,
(	9810	)	,
(	9809	)	,
(	9807	)	,
(	9806	)	,
(	9804	)	,
(	9802	)	,
(	9801	)	,
(	9799	)	,
(	9797	)	,
(	9796	)	,
(	9794	)	,
(	9793	)	,
(	9791	)	,
(	9789	)	,
(	9788	)	,
(	9786	)	,
(	9785	)	,
(	9783	)	,
(	9781	)	,
(	9780	)	,
(	9778	)	,
(	9776	)	,
(	9775	)	,
(	9773	)	,
(	9772	)	,
(	9770	)	,
(	9768	)	,
(	9767	)	,
(	9765	)	,
(	9763	)	,
(	9762	)	,
(	9760	)	,
(	9759	)	,
(	9757	)	,
(	9755	)	,
(	9754	)	,
(	9752	)	,
(	9751	)	,
(	9749	)	,
(	9747	)	,
(	9746	)	,
(	9744	)	,
(	9742	)	,
(	9741	)	,
(	9739	)	,
(	9738	)	,
(	9736	)	,
(	9734	)	,
(	9733	)	,
(	9731	)	,
(	9729	)	,
(	9728	)	,
(	9726	)	,
(	9725	)	,
(	9723	)	,
(	9721	)	,
(	9720	)	,
(	9718	)	,
(	9716	)	,
(	9715	)	,
(	9713	)	,
(	9712	)	,
(	9710	)	,
(	9708	)	,
(	9707	)	,
(	9705	)	,
(	9704	)	,
(	9702	)	,
(	9700	)	,
(	9699	)	,
(	9697	)	,
(	9695	)	,
(	9694	)	,
(	9692	)	,
(	9691	)	,
(	9689	)	,
(	9687	)	,
(	9686	)	,
(	9684	)	,
(	9682	)	,
(	9681	)	,
(	9679	)	,
(	9678	)	,
(	9676	)	,
(	9674	)	,
(	9673	)	,
(	9671	)	,
(	9670	)	,
(	9668	)	,
(	9666	)	,
(	9665	)	,
(	9663	)	,
(	9661	)	,
(	9660	)	,
(	9658	)	,
(	9657	)	,
(	9655	)	,
(	9653	)	,
(	9652	)	,
(	9650	)	,
(	9648	)	,
(	9647	)	,
(	9645	)	,
(	9644	)	,
(	9642	)	,
(	9640	)	,
(	9639	)	,
(	9637	)	,
(	9635	)	,
(	9634	)	,
(	9632	)	,
(	9631	)	,
(	9629	)	,
(	9627	)	,
(	9626	)	,
(	9624	)	,
(	9623	)	,
(	9621	)	,
(	9619	)	,
(	9618	)	,
(	9616	)	,
(	9614	)	,
(	9613	)	,
(	9611	)	,
(	9610	)	,
(	9608	)	,
(	9606	)	,
(	9605	)	,
(	9603	)	,
(	9601	)	,
(	9600	)	,
(	9598	)	,
(	9597	)	,
(	9595	)	,
(	9593	)	,
(	9592	)	,
(	9590	)	,
(	9589	)	,
(	9587	)	,
(	9585	)	,
(	9584	)	,
(	9582	)	,
(	9580	)	,
(	9579	)	,
(	9577	)	,
(	9576	)	,
(	9574	)	,
(	9572	)	,
(	9571	)	,
(	9569	)	,
(	9567	)	,
(	9566	)	,
(	9564	)	,
(	9563	)	,
(	9561	)	,
(	9559	)	,
(	9558	)	,
(	9556	)	,
(	9554	)	,
(	9553	)	,
(	9551	)	,
(	9550	)	,
(	9548	)	,
(	9546	)	,
(	9545	)	,
(	9543	)	,
(	9542	)	,
(	9540	)	,
(	9538	)	,
(	9537	)	,
(	9535	)	,
(	9533	)	,
(	9532	)	,
(	9530	)	,
(	9529	)	,
(	9527	)	,
(	9525	)	,
(	9524	)	,
(	9522	)	,
(	9520	)	,
(	9519	)	,
(	9517	)	,
(	9516	)	,
(	9514	)	,
(	9512	)	,
(	9511	)	,
(	9509	)	,
(	9508	)	,
(	9506	)	,
(	9504	)	,
(	9503	)	,
(	9501	)	,
(	9499	)	,
(	9498	)	,
(	9496	)	,
(	9495	)	,
(	9493	)	,
(	9491	)	,
(	9490	)	,
(	9488	)	,
(	9486	)	,
(	9485	)	,
(	9483	)	,
(	9482	)	,
(	9480	)	,
(	9478	)	,
(	9477	)	,
(	9475	)	,
(	9473	)	,
(	9472	)	,
(	9470	)	,
(	9469	)	,
(	9467	)	,
(	9465	)	,
(	9464	)	,
(	9462	)	,
(	9461	)	,
(	9459	)	,
(	9457	)	,
(	9456	)	,
(	9454	)	,
(	9452	)	,
(	9451	)	,
(	9449	)	,
(	9448	)	,
(	9446	)	,
(	9444	)	,
(	9443	)	,
(	9441	)	,
(	9439	)	,
(	9438	)	,
(	9436	)	,
(	9435	)	,
(	9433	)	,
(	9431	)	,
(	9430	)	,
(	9428	)	,
(	9427	)	,
(	9425	)	,
(	9423	)	,
(	9422	)	,
(	9420	)	,
(	9418	)	,
(	9417	)	,
(	9415	)	,
(	9414	)	,
(	9412	)	,
(	9410	)	,
(	9409	)	,
(	9407	)	,
(	9405	)	,
(	9404	)	,
(	9402	)	,
(	9401	)	,
(	9399	)	,
(	9397	)	,
(	9396	)	,
(	9394	)	,
(	9392	)	,
(	9391	)	,
(	9389	)	,
(	9388	)	,
(	9386	)	,
(	9384	)	,
(	9383	)	,
(	9381	)	,
(	9380	)	,
(	9378	)	,
(	9376	)	,
(	9375	)	,
(	9373	)	,
(	9371	)	,
(	9370	)	,
(	9368	)	,
(	9367	)	,
(	9365	)	,
(	9363	)	,
(	9362	)	,
(	9360	)	,
(	9358	)	,
(	9357	)	,
(	9355	)	,
(	9354	)	,
(	9352	)	,
(	9350	)	,
(	9349	)	,
(	9347	)	,
(	9346	)	,
(	9344	)	,
(	9342	)	,
(	9341	)	,
(	9339	)	,
(	9337	)	,
(	9336	)	,
(	9334	)	,
(	9333	)	,
(	9331	)	,
(	9329	)	,
(	9328	)	,
(	9326	)	,
(	9324	)	,
(	9323	)	,
(	9321	)	,
(	9320	)	,
(	9318	)	,
(	9316	)	,
(	9315	)	,
(	9313	)	,
(	9311	)	,
(	9310	)	,
(	9308	)	,
(	9307	)	,
(	9305	)	,
(	9303	)	,
(	9302	)	,
(	9300	)	,
(	9299	)	,
(	9297	)	,
(	9295	)	,
(	9294	)	,
(	9292	)	,
(	9290	)	,
(	9289	)	,
(	9287	)	,
(	9286	)	,
(	9284	)	,
(	9282	)	,
(	9281	)	,
(	9279	)	,
(	9277	)	,
(	9276	)	,
(	9274	)	,
(	9273	)	,
(	9271	)	,
(	9269	)	,
(	9268	)	,
(	9266	)	,
(	9265	)	,
(	9263	)	,
(	9261	)	,
(	9260	)	,
(	9258	)	,
(	9256	)	,
(	9255	)	,
(	9253	)	,
(	9252	)	,
(	9250	)	,
(	9248	)	,
(	9247	)	,
(	9245	)	,
(	9243	)	,
(	9242	)	,
(	9240	)	,
(	9239	)	,
(	9237	)	,
(	9235	)	,
(	9234	)	,
(	9232	)	,
(	9230	)	,
(	9229	)	,
(	9227	)	,
(	9226	)	,
(	9224	)	,
(	9222	)	,
(	9221	)	,
(	9219	)	,
(	9218	)	,
(	9216	)	,
(	9214	)	,
(	9213	)	,
(	9211	)	,
(	9209	)	,
(	9208	)	,
(	9206	)	,
(	9205	)	,
(	9203	)	,
(	9201	)	,
(	9200	)	,
(	9198	)	,
(	9196	)	,
(	9195	)	,
(	9193	)	,
(	9192	)	,
(	9190	)	,
(	9188	)	,
(	9187	)	,
(	9185	)	,
(	9184	)	,
(	9182	)	,
(	9180	)	,
(	9179	)	,
(	9177	)	,
(	9175	)	,
(	9174	)	,
(	9172	)	,
(	9171	)	,
(	9169	)	,
(	9167	)	,
(	9166	)	,
(	9164	)	,
(	9162	)	,
(	9161	)	,
(	9159	)	,
(	9158	)	,
(	9156	)	,
(	9154	)	,
(	9153	)	,
(	9151	)	,
(	9149	)	,
(	9148	)	,
(	9146	)	,
(	9145	)	,
(	9143	)	,
(	9141	)	,
(	9140	)	,
(	9138	)	,
(	9137	)	,
(	9135	)	,
(	9133	)	,
(	9132	)	,
(	9130	)	,
(	9128	)	,
(	9127	)	,
(	9125	)	,
(	9124	)	,
(	9122	)	,
(	9120	)	,
(	9119	)	,
(	9117	)	,
(	9115	)	,
(	9114	)	,
(	9112	)	,
(	9111	)	,
(	9109	)	,
(	9107	)	,
(	9106	)	,
(	9104	)	,
(	9103	)	,
(	9101	)	,
(	9099	)	,
(	9098	)	,
(	9096	)	,
(	9094	)	,
(	9093	)	,
(	9091	)	,
(	9090	)	,
(	9088	)	,
(	9086	)	,
(	9085	)	,
(	9083	)	,
(	9081	)	,
(	9080	)	,
(	9078	)	,
(	9077	)	,
(	9075	)	,
(	9073	)	,
(	9072	)	,
(	9070	)	,
(	9068	)	,
(	9067	)	,
(	9065	)	,
(	9064	)	,
(	9062	)	,
(	9060	)	,
(	9059	)	,
(	9057	)	,
(	9056	)	,
(	9054	)	,
(	9052	)	,
(	9051	)	,
(	9049	)	,
(	9047	)	,
(	9046	)	,
(	9044	)	,
(	9043	)	,
(	9041	)	,
(	9039	)	,
(	9038	)	,
(	9036	)	,
(	9034	)	,
(	9033	)	,
(	9031	)	,
(	9030	)	,
(	9028	)	,
(	9026	)	,
(	9025	)	,
(	9023	)	,
(	9022	)	,
(	9020	)	,
(	9018	)	,
(	9017	)	,
(	9015	)	,
(	9013	)	,
(	9012	)	,
(	9010	)	,
(	9009	)	,
(	9007	)	,
(	9005	)	,
(	9004	)	,
(	9002	)	,
(	9000	)	,
(	8999	)	,
(	8997	)	,
(	8996	)	,
(	8994	)	,
(	8992	)	,
(	8991	)	,
(	8989	)	,
(	8987	)	,
(	8986	)	,
(	8984	)	,
(	8983	)	,
(	8981	)	,
(	8979	)	,
(	8978	)	,
(	8976	)	,
(	8975	)	,
(	8973	)	,
(	8971	)	,
(	8970	)	,
(	8968	)	,
(	8966	)	,
(	8965	)	,
(	8963	)	,
(	8962	)	,
(	8960	)	,
(	8958	)	,
(	8957	)	,
(	8955	)	,
(	8953	)	,
(	8952	)	,
(	8950	)	,
(	8949	)	,
(	8947	)	,
(	8945	)	,
(	8944	)	,
(	8942	)	,
(	8941	)	,
(	8939	)	,
(	8937	)	,
(	8936	)	,
(	8934	)	,
(	8932	)	,
(	8931	)	,
(	8929	)	,
(	8928	)	,
(	8926	)	,
(	8924	)	,
(	8923	)	,
(	8921	)	,
(	8919	)	,
(	8918	)	,
(	8916	)	,
(	8915	)	,
(	8913	)	,
(	8911	)	,
(	8910	)	,
(	8908	)	,
(	8906	)	,
(	8905	)	,
(	8903	)	,
(	8902	)	,
(	8900	)	,
(	8898	)	,
(	8897	)	,
(	8895	)	,
(	8894	)	,
(	8892	)	,
(	8890	)	,
(	8889	)	,
(	8887	)	,
(	8885	)	,
(	8884	)	,
(	8882	)	,
(	8881	)	,
(	8879	)	,
(	8877	)	,
(	8876	)	,
(	8874	)	,
(	8872	)	,
(	8871	)	,
(	8869	)	,
(	8868	)	,
(	8866	)	,
(	8864	)	,
(	8863	)	,
(	8861	)	,
(	8860	)	,
(	8858	)	,
(	8856	)	,
(	8855	)	,
(	8853	)	,
(	8851	)	,
(	8850	)	,
(	8848	)	,
(	8847	)	,
(	8845	)	,
(	8843	)	,
(	8842	)	,
(	8840	)	,
(	8838	)	,
(	8837	)	,
(	8835	)	,
(	8834	)	,
(	8832	)	,
(	8830	)	,
(	8829	)	,
(	8827	)	,
(	8825	)	,
(	8824	)	,
(	8822	)	,
(	8821	)	,
(	8819	)	,
(	8817	)	,
(	8816	)	,
(	8814	)	,
(	8813	)	,
(	8811	)	,
(	8809	)	,
(	8808	)	,
(	8806	)	,
(	8804	)	,
(	8803	)	,
(	8801	)	,
(	8800	)	,
(	8798	)	,
(	8796	)	,
(	8795	)	,
(	8793	)	,
(	8791	)	,
(	8790	)	,
(	8788	)	,
(	8787	)	,
(	8785	)	,
(	8783	)	,
(	8782	)	,
(	8780	)	,
(	8779	)	,
(	8777	)	,
(	8775	)	,
(	8774	)	,
(	8772	)	,
(	8770	)	,
(	8769	)	,
(	8767	)	,
(	8766	)	,
(	8764	)	,
(	8762	)	,
(	8761	)	,
(	8759	)	,
(	8757	)	,
(	8756	)	,
(	8754	)	,
(	8753	)	,
(	8751	)	,
(	8749	)	,
(	8748	)	,
(	8746	)	,
(	8744	)	,
(	8743	)	,
(	8741	)	,
(	8740	)	,
(	8738	)	,
(	8736	)	,
(	8735	)	,
(	8733	)	,
(	8732	)	,
(	8730	)	,
(	8728	)	,
(	8727	)	,
(	8725	)	,
(	8723	)	,
(	8722	)	,
(	8720	)	,
(	8719	)	,
(	8717	)	,
(	8715	)	,
(	8714	)	,
(	8712	)	,
(	8710	)	,
(	8709	)	,
(	8707	)	,
(	8706	)	,
(	8704	)	,
(	8702	)	,
(	8701	)	,
(	8699	)	,
(	8698	)	,
(	8696	)	,
(	8694	)	,
(	8693	)	,
(	8691	)	,
(	8689	)	,
(	8688	)	,
(	8686	)	,
(	8685	)	,
(	8683	)	,
(	8681	)	,
(	8680	)	,
(	8678	)	,
(	8676	)	,
(	8675	)	,
(	8673	)	,
(	8672	)	,
(	8670	)	,
(	8668	)	,
(	8667	)	,
(	8665	)	,
(	8663	)	,
(	8662	)	,
(	8660	)	,
(	8659	)	,
(	8657	)	,
(	8655	)	,
(	8654	)	,
(	8652	)	,
(	8651	)	,
(	8649	)	,
(	8647	)	,
(	8646	)	,
(	8644	)	,
(	8642	)	,
(	8641	)	,
(	8639	)	,
(	8638	)	,
(	8636	)	,
(	8634	)	,
(	8633	)	,
(	8631	)	,
(	8629	)	,
(	8628	)	,
(	8626	)	,
(	8625	)	,
(	8623	)	,
(	8621	)	,
(	8620	)	,
(	8618	)	,
(	8617	)	,
(	8615	)	,
(	8613	)	,
(	8612	)	,
(	8610	)	,
(	8608	)	,
(	8607	)	,
(	8605	)	,
(	8604	)	,
(	8602	)	,
(	8600	)	,
(	8599	)	,
(	8597	)	,
(	8595	)	,
(	8594	)	,
(	8592	)	,
(	8591	)	,
(	8589	)	,
(	8587	)	,
(	8586	)	,
(	8584	)	,
(	8582	)	,
(	8581	)	,
(	8579	)	,
(	8578	)	,
(	8576	)	,
(	8574	)	,
(	8573	)	,
(	8571	)	,
(	8570	)	,
(	8568	)	,
(	8566	)	,
(	8565	)	,
(	8563	)	,
(	8561	)	,
(	8560	)	,
(	8558	)	,
(	8557	)	,
(	8555	)	,
(	8553	)	,
(	8552	)	,
(	8550	)	,
(	8548	)	,
(	8547	)	,
(	8545	)	,
(	8544	)	,
(	8542	)	,
(	8540	)	,
(	8539	)	,
(	8537	)	,
(	8536	)	,
(	8534	)	,
(	8532	)	,
(	8531	)	,
(	8529	)	,
(	8527	)	,
(	8526	)	,
(	8524	)	,
(	8523	)	,
(	8521	)	,
(	8519	)	,
(	8518	)	,
(	8516	)	,
(	8514	)	,
(	8513	)	,
(	8511	)	,
(	8510	)	,
(	8508	)	,
(	8506	)	,
(	8505	)	,
(	8503	)	,
(	8501	)	,
(	8500	)	,
(	8498	)	,
(	8497	)	,
(	8495	)	,
(	8493	)	,
(	8492	)	,
(	8490	)	,
(	8489	)	,
(	8487	)	,
(	8485	)	,
(	8484	)	,
(	8482	)	,
(	8480	)	,
(	8479	)	,
(	8477	)	,
(	8476	)	,
(	8474	)	,
(	8472	)	,
(	8471	)	,
(	8469	)	,
(	8467	)	,
(	8466	)	,
(	8464	)	,
(	8463	)	,
(	8461	)	,
(	8459	)	,
(	8458	)	,
(	8456	)	,
(	8455	)	,
(	8453	)	,
(	8451	)	,
(	8450	)	,
(	8448	)	,
(	8446	)	,
(	8445	)	,
(	8443	)	,
(	8442	)	,
(	8440	)	,
(	8438	)	,
(	8437	)	,
(	8435	)	,
(	8433	)	,
(	8432	)	,
(	8430	)	,
(	8429	)	,
(	8427	)	,
(	8425	)	,
(	8424	)	,
(	8422	)	,
(	8420	)	,
(	8419	)	,
(	8417	)	,
(	8416	)	,
(	8414	)	,
(	8412	)	,
(	8411	)	,
(	8409	)	,
(	8408	)	,
(	8406	)	,
(	8404	)	,
(	8403	)	,
(	8401	)	,
(	8399	)	,
(	8398	)	,
(	8396	)	,
(	8395	)	,
(	8393	)	,
(	8391	)	,
(	8390	)	,
(	8388	)	,
(	8386	)	,
(	8385	)	,
(	8383	)	,
(	8382	)	,
(	8380	)	,
(	8378	)	,
(	8377	)	,
(	8375	)	,
(	8374	)	,
(	8372	)	,
(	8370	)	,
(	8369	)	,
(	8367	)	,
(	8365	)	,
(	8364	)	,
(	8362	)	,
(	8361	)	,
(	8359	)	,
(	8357	)	,
(	8356	)	,
(	8354	)	,
(	8352	)	,
(	8351	)	,
(	8349	)	,
(	8348	)	,
(	8346	)	,
(	8344	)	,
(	8343	)	,
(	8341	)	,
(	8339	)	,
(	8338	)	,
(	8336	)	,
(	8335	)	,
(	8333	)	,
(	8331	)	,
(	8330	)	,
(	8328	)	,
(	8327	)	,
(	8325	)	,
(	8323	)	,
(	8322	)	,
(	8320	)	,
(	8318	)	,
(	8317	)	,
(	8315	)	,
(	8314	)	,
(	8312	)	,
(	8310	)	,
(	8309	)	,
(	8307	)	,
(	8305	)	,
(	8304	)	,
(	8302	)	,
(	8301	)	,
(	8299	)	,
(	8297	)	,
(	8296	)	,
(	8294	)	,
(	8293	)	,
(	8291	)	,
(	8289	)	,
(	8288	)	,
(	8286	)	,
(	8284	)	,
(	8283	)	,
(	8281	)	,
(	8280	)	,
(	8278	)	,
(	8276	)	,
(	8275	)	,
(	8273	)	,
(	8271	)	,
(	8270	)	,
(	8268	)	,
(	8267	)	,
(	8265	)	,
(	8263	)	,
(	8262	)	,
(	8260	)	,
(	8258	)	,
(	8257	)	,
(	8255	)	,
(	8254	)	,
(	8252	)	,
(	8250	)	,
(	8249	)	,
(	8247	)	,
(	8246	)	,
(	8244	)	,
(	8242	)	,
(	8241	)	,
(	8239	)	,
(	8237	)	,
(	8236	)	,
(	8234	)	,
(	8233	)	,
(	8231	)	,
(	8229	)	,
(	8228	)	,
(	8226	)	,
(	8224	)	,
(	8223	)	,
(	8221	)	,
(	8220	)	,
(	8218	)	,
(	8216	)	,
(	8215	)	,
(	8213	)	,
(	8212	)	,
(	8210	)	,
(	8208	)	,
(	8207	)	,
(	8205	)	,
(	8203	)	,
(	8202	)	,
(	8200	)	,
(	8199	)	,
(	8197	)	,
(	8195	)	,
(	8194	)	,
(	8192	)	,
(	8190	)	,
(	8189	)	,
(	8187	)	,
(	8186	)	,
(	8184	)	,
(	8182	)	,
(	8181	)	,
(	8179	)	,
(	8177	)	,
(	8176	)	,
(	8174	)	,
(	8173	)	,
(	8171	)	,
(	8169	)	,
(	8168	)	,
(	8166	)	,
(	8165	)	,
(	8163	)	,
(	8161	)	,
(	8160	)	,
(	8158	)	,
(	8156	)	,
(	8155	)	,
(	8153	)	,
(	8152	)	,
(	8150	)	,
(	8148	)	,
(	8147	)	,
(	8145	)	,
(	8143	)	,
(	8142	)	,
(	8140	)	,
(	8139	)	,
(	8137	)	,
(	8135	)	,
(	8134	)	,
(	8132	)	,
(	8131	)	,
(	8129	)	,
(	8127	)	,
(	8126	)	,
(	8124	)	,
(	8122	)	,
(	8121	)	,
(	8119	)	,
(	8118	)	,
(	8116	)	,
(	8114	)	,
(	8113	)	,
(	8111	)	,
(	8109	)	,
(	8108	)	,
(	8106	)	,
(	8105	)	,
(	8103	)	,
(	8101	)	,
(	8100	)	,
(	8098	)	,
(	8096	)	,
(	8095	)	,
(	8093	)	,
(	8092	)	,
(	8090	)	,
(	8088	)	,
(	8087	)	,
(	8085	)	,
(	8084	)	,
(	8082	)	,
(	8080	)	,
(	8079	)	,
(	8077	)	,
(	8075	)	,
(	8074	)	,
(	8072	)	,
(	8071	)	,
(	8069	)	,
(	8067	)	,
(	8066	)	,
(	8064	)	,
(	8062	)	,
(	8061	)	,
(	8059	)	,
(	8058	)	,
(	8056	)	,
(	8054	)	,
(	8053	)	,
(	8051	)	,
(	8050	)	,
(	8048	)	,
(	8046	)	,
(	8045	)	,
(	8043	)	,
(	8041	)	,
(	8040	)	,
(	8038	)	,
(	8037	)	,
(	8035	)	,
(	8033	)	,
(	8032	)	,
(	8030	)	,
(	8028	)	,
(	8027	)	,
(	8025	)	,
(	8024	)	,
(	8022	)	,
(	8020	)	,
(	8019	)	,
(	8017	)	,
(	8015	)	,
(	8014	)	,
(	8012	)	,
(	8011	)	,
(	8009	)	,
(	8007	)	,
(	8006	)	,
(	8004	)	,
(	8003	)	,
(	8001	)	,
(	7999	)	,
(	7998	)	,
(	7996	)	,
(	7994	)	,
(	7993	)	,
(	7991	)	,
(	7990	)	,
(	7988	)	,
(	7986	)	,
(	7985	)	,
(	7983	)	,
(	7981	)	,
(	7980	)	,
(	7978	)	,
(	7977	)	,
(	7975	)	,
(	7973	)	,
(	7972	)	,
(	7970	)	,
(	7969	)	,
(	7967	)	,
(	7965	)	,
(	7964	)	,
(	7962	)	,
(	7960	)	,
(	7959	)	,
(	7957	)	,
(	7956	)	,
(	7954	)	,
(	7952	)	,
(	7951	)	,
(	7949	)	,
(	7947	)	,
(	7946	)	,
(	7944	)	,
(	7943	)	,
(	7941	)	,
(	7939	)	,
(	7938	)	,
(	7936	)	,
(	7934	)	,
(	7933	)	,
(	7931	)	,
(	7930	)	,
(	7928	)	,
(	7926	)	,
(	7925	)	,
(	7923	)	,
(	7922	)	,
(	7920	)	,
(	7918	)	,
(	7917	)	,
(	7915	)	,
(	7913	)	,
(	7912	)	,
(	7910	)	,
(	7909	)	,
(	7907	)	,
(	7905	)	,
(	7904	)	,
(	7902	)	,
(	7900	)	,
(	7899	)	,
(	7897	)	,
(	7896	)	,
(	7894	)	,
(	7892	)	,
(	7891	)	,
(	7889	)	,
(	7888	)	,
(	7886	)	,
(	7884	)	,
(	7883	)	,
(	7881	)	,
(	7879	)	,
(	7878	)	,
(	7876	)	,
(	7875	)	,
(	7873	)	,
(	7871	)	,
(	7870	)	,
(	7868	)	,
(	7866	)	,
(	7865	)	,
(	7863	)	,
(	7862	)	,
(	7860	)	,
(	7858	)	,
(	7857	)	,
(	7855	)	,
(	7853	)	,
(	7852	)	,
(	7850	)	,
(	7849	)	,
(	7847	)	,
(	7845	)	,
(	7844	)	,
(	7842	)	,
(	7841	)	,
(	7839	)	,
(	7837	)	,
(	7836	)	,
(	7834	)	,
(	7832	)	,
(	7831	)	,
(	7829	)	,
(	7828	)	,
(	7826	)	,
(	7824	)	,
(	7823	)	,
(	7821	)	,
(	7819	)	,
(	7818	)	,
(	7816	)	,
(	7815	)	,
(	7813	)	,
(	7811	)	,
(	7810	)	,
(	7808	)	,
(	7807	)	,
(	7805	)	,
(	7803	)	,
(	7802	)	,
(	7800	)	,
(	7798	)	,
(	7797	)	,
(	7795	)	,
(	7794	)	,
(	7792	)	,
(	7790	)	,
(	7789	)	,
(	7787	)	,
(	7785	)	,
(	7784	)	,
(	7782	)	,
(	7781	)	,
(	7779	)	,
(	7777	)	,
(	7776	)	,
(	7774	)	,
(	7772	)	,
(	7771	)	,
(	7769	)	,
(	7768	)	,
(	7766	)	,
(	7764	)	,
(	7763	)	,
(	7761	)	,
(	7760	)	,
(	7758	)	,
(	7756	)	,
(	7755	)	,
(	7753	)	,
(	7751	)	,
(	7750	)	,
(	7748	)	,
(	7747	)	,
(	7745	)	,
(	7743	)	,
(	7742	)	,
(	7740	)	,
(	7738	)	,
(	7737	)	,
(	7735	)	,
(	7734	)	,
(	7732	)	,
(	7730	)	,
(	7729	)	,
(	7727	)	,
(	7726	)	,
(	7724	)	,
(	7722	)	,
(	7721	)	,
(	7719	)	,
(	7717	)	,
(	7716	)	,
(	7714	)	,
(	7713	)	,
(	7711	)	,
(	7709	)	,
(	7708	)	,
(	7706	)	,
(	7704	)	,
(	7703	)	,
(	7701	)	,
(	7700	)	,
(	7698	)	,
(	7696	)	,
(	7695	)	,
(	7693	)	,
(	7691	)	,
(	7690	)	,
(	7688	)	,
(	7687	)	,
(	7685	)	,
(	7683	)	,
(	7682	)	,
(	7680	)	,
(	7679	)	,
(	7677	)	,
(	7675	)	,
(	7674	)	,
(	7672	)	,
(	7670	)	,
(	7669	)	,
(	7667	)	,
(	7666	)	,
(	7664	)	,
(	7662	)	,
(	7661	)	,
(	7659	)	,
(	7657	)	,
(	7656	)	,
(	7654	)	,
(	7653	)	,
(	7651	)	,
(	7649	)	,
(	7648	)	,
(	7646	)	,
(	7645	)	,
(	7643	)	,
(	7641	)	,
(	7640	)	,
(	7638	)	,
(	7636	)	,
(	7635	)	,
(	7633	)	,
(	7632	)	,
(	7630	)	,
(	7628	)	,
(	7627	)	,
(	7625	)	,
(	7623	)	,
(	7622	)	,
(	7620	)	,
(	7619	)	,
(	7617	)	,
(	7615	)	,
(	7614	)	,
(	7612	)	,
(	7610	)	,
(	7609	)	,
(	7607	)	,
(	7606	)	,
(	7604	)	,
(	7602	)	,
(	7601	)	,
(	7599	)	,
(	7598	)	,
(	7596	)	,
(	7594	)	,
(	7593	)	,
(	7591	)	,
(	7589	)	,
(	7588	)	,
(	7586	)	,
(	7585	)	,
(	7583	)	,
(	7581	)	,
(	7580	)	,
(	7578	)	,
(	7576	)	,
(	7575	)	,
(	7573	)	,
(	7572	)	,
(	7570	)	,
(	7568	)	,
(	7567	)	,
(	7565	)	,
(	7564	)	,
(	7562	)	,
(	7560	)	,
(	7559	)	,
(	7557	)	,
(	7555	)	,
(	7554	)	,
(	7552	)	,
(	7551	)	,
(	7549	)	,
(	7547	)	,
(	7546	)	,
(	7544	)	,
(	7542	)	,
(	7541	)	,
(	7539	)	,
(	7538	)	,
(	7536	)	,
(	7534	)	,
(	7533	)	,
(	7531	)	,
(	7529	)	,
(	7528	)	,
(	7526	)	,
(	7525	)	,
(	7523	)	,
(	7521	)	,
(	7520	)	,
(	7518	)	,
(	7517	)	,
(	7515	)	,
(	7513	)	,
(	7512	)	,
(	7510	)	,
(	7508	)	,
(	7507	)	,
(	7505	)	,
(	7504	)	,
(	7502	)	,
(	7500	)	,
(	7499	)	,
(	7497	)	,
(	7495	)	,
(	7494	)	,
(	7492	)	,
(	7491	)	,
(	7489	)	,
(	7487	)	,
(	7486	)	,
(	7484	)	,
(	7483	)	,
(	7481	)	,
(	7479	)	,
(	7478	)	,
(	7476	)	,
(	7474	)	,
(	7473	)	,
(	7471	)	,
(	7470	)	,
(	7468	)	,
(	7466	)	,
(	7465	)	,
(	7463	)	,
(	7461	)	,
(	7460	)	,
(	7458	)	,
(	7457	)	,
(	7455	)	,
(	7453	)	,
(	7452	)	,
(	7450	)	,
(	7448	)	,
(	7447	)	,
(	7445	)	,
(	7444	)	,
(	7442	)	,
(	7440	)	,
(	7439	)	,
(	7437	)	,
(	7436	)	,
(	7434	)	,
(	7432	)	,
(	7431	)	,
(	7429	)	,
(	7427	)	,
(	7426	)	,
(	7424	)	,
(	7423	)	,
(	7421	)	,
(	7419	)	,
(	7418	)	,
(	7416	)	,
(	7414	)	,
(	7413	)	,
(	7411	)	,
(	7410	)	,
(	7408	)	,
(	7406	)	,
(	7405	)	,
(	7403	)	,
(	7402	)	,
(	7400	)	,
(	7398	)	,
(	7397	)	,
(	7395	)	,
(	7393	)	,
(	7392	)	,
(	7390	)	,
(	7389	)	,
(	7387	)	,
(	7385	)	,
(	7384	)	,
(	7382	)	,
(	7380	)	,
(	7379	)	,
(	7377	)	,
(	7376	)	,
(	7374	)	,
(	7372	)	,
(	7371	)	,
(	7369	)	,
(	7367	)	,
(	7366	)	,
(	7364	)	,
(	7363	)	,
(	7361	)	,
(	7359	)	,
(	7358	)	,
(	7356	)	,
(	7355	)	,
(	7353	)	,
(	7351	)	,
(	7350	)	,
(	7348	)	,
(	7346	)	,
(	7345	)	,
(	7343	)	,
(	7342	)	,
(	7340	)	,
(	7338	)	,
(	7337	)	,
(	7335	)	,
(	7333	)	,
(	7332	)	,
(	7330	)	,
(	7329	)	,
(	7327	)	,
(	7325	)	,
(	7324	)	,
(	7322	)	,
(	7321	)	,
(	7319	)	,
(	7317	)	,
(	7316	)	,
(	7314	)	,
(	7312	)	,
(	7311	)	,
(	7309	)	,
(	7308	)	,
(	7306	)	,
(	7304	)	,
(	7303	)	,
(	7301	)	,
(	7299	)	,
(	7298	)	,
(	7296	)	,
(	7295	)	,
(	7293	)	,
(	7291	)	,
(	7290	)	,
(	7288	)	,
(	7286	)	,
(	7285	)	,
(	7283	)	,
(	7282	)	,
(	7280	)	,
(	7278	)	,
(	7277	)	,
(	7275	)	,
(	7274	)	,
(	7272	)	,
(	7270	)	,
(	7269	)	,
(	7267	)	,
(	7265	)	,
(	7264	)	,
(	7262	)	,
(	7261	)	,
(	7259	)	,
(	7257	)	,
(	7256	)	,
(	7254	)	,
(	7252	)	,
(	7251	)	,
(	7249	)	,
(	7248	)	,
(	7246	)	,
(	7244	)	,
(	7243	)	,
(	7241	)	,
(	7240	)	,
(	7238	)	,
(	7236	)	,
(	7235	)	,
(	7233	)	,
(	7231	)	,
(	7230	)	,
(	7228	)	,
(	7227	)	,
(	7225	)	,
(	7223	)	,
(	7222	)	,
(	7220	)	,
(	7218	)	,
(	7217	)	,
(	7215	)	,
(	7214	)	,
(	7212	)	,
(	7210	)	,
(	7209	)	,
(	7207	)	,
(	7205	)	,
(	7204	)	,
(	7202	)	,
(	7201	)	,
(	7199	)	,
(	7197	)	,
(	7196	)	,
(	7194	)	,
(	7193	)	,
(	7191	)	,
(	7189	)	,
(	7188	)	,
(	7186	)	,
(	7184	)	,
(	7183	)	,
(	7181	)	,
(	7180	)	,
(	7178	)	,
(	7176	)	,
(	7175	)	,
(	7173	)	,
(	7171	)	,
(	7170	)	,
(	7168	)	,
(	7167	)	,
(	7165	)	,
(	7163	)	,
(	7162	)	,
(	7160	)	,
(	7159	)	,
(	7157	)	,
(	7155	)	,
(	7154	)	,
(	7152	)	,
(	7150	)	,
(	7149	)	,
(	7147	)	,
(	7146	)	,
(	7144	)	,
(	7142	)	,
(	7141	)	,
(	7139	)	,
(	7137	)	,
(	7136	)	,
(	7134	)	,
(	7133	)	,
(	7131	)	,
(	7129	)	,
(	7128	)	,
(	7126	)	,
(	7124	)	,
(	7123	)	,
(	7121	)	,
(	7120	)	,
(	7118	)	,
(	7116	)	,
(	7115	)	,
(	7113	)	,
(	7112	)	,
(	7110	)	,
(	7108	)	,
(	7107	)	,
(	7105	)	,
(	7103	)	,
(	7102	)	,
(	7100	)	,
(	7099	)	,
(	7097	)	,
(	7095	)	,
(	7094	)	,
(	7092	)	,
(	7090	)	,
(	7089	)	,
(	7087	)	,
(	7086	)	,
(	7084	)	,
(	7082	)	,
(	7081	)	,
(	7079	)	,
(	7078	)	,
(	7076	)	,
(	7074	)	,
(	7073	)	,
(	7071	)	,
(	7069	)	,
(	7068	)	,
(	7066	)	,
(	7065	)	,
(	7063	)	,
(	7061	)	,
(	7060	)	,
(	7058	)	,
(	7056	)	,
(	7055	)	,
(	7053	)	,
(	7052	)	,
(	7050	)	,
(	7048	)	,
(	7047	)	,
(	7045	)	,
(	7043	)	,
(	7042	)	,
(	7040	)	,
(	7039	)	,
(	7037	)	,
(	7035	)	,
(	7034	)	,
(	7032	)	,
(	7031	)	,
(	7029	)	,
(	7027	)	,
(	7026	)	,
(	7024	)	,
(	7022	)	,
(	7021	)	,
(	7019	)	,
(	7018	)	,
(	7016	)	,
(	7014	)	,
(	7013	)	,
(	7011	)	,
(	7009	)	,
(	7008	)	,
(	7006	)	,
(	7005	)	,
(	7003	)	,
(	7001	)	,
(	7000	)	,
(	6998	)	,
(	6997	)	,
(	6995	)	,
(	6993	)	,
(	6992	)	,
(	6990	)	,
(	6988	)	,
(	6987	)	,
(	6985	)	,
(	6984	)	,
(	6982	)	,
(	6980	)	,
(	6979	)	,
(	6977	)	,
(	6975	)	,
(	6974	)	,
(	6972	)	,
(	6971	)	,
(	6969	)	,
(	6967	)	,
(	6966	)	,
(	6964	)	,
(	6962	)	,
(	6961	)	,
(	6959	)	,
(	6958	)	,
(	6956	)	,
(	6954	)	,
(	6953	)	,
(	6951	)	,
(	6950	)	,
(	6948	)	,
(	6946	)	,
(	6945	)	,
(	6943	)	,
(	6941	)	,
(	6940	)	,
(	6938	)	,
(	6937	)	,
(	6935	)	,
(	6933	)	,
(	6932	)	,
(	6930	)	,
(	6928	)	,
(	6927	)	,
(	6925	)	,
(	6924	)	,
(	6922	)	,
(	6920	)	,
(	6919	)	,
(	6917	)	,
(	6916	)	,
(	6914	)	,
(	6912	)	,
(	6911	)	,
(	6909	)	,
(	6907	)	,
(	6906	)	,
(	6904	)	,
(	6903	)	,
(	6901	)	,
(	6899	)	,
(	6898	)	,
(	6896	)	,
(	6894	)	,
(	6893	)	,
(	6891	)	,
(	6890	)	,
(	6888	)	,
(	6886	)	,
(	6885	)	,
(	6883	)	,
(	6881	)	,
(	6880	)	,
(	6878	)	,
(	6877	)	,
(	6875	)	,
(	6873	)	,
(	6872	)	,
(	6870	)	,
(	6869	)	,
(	6867	)	,
(	6865	)	,
(	6864	)	,
(	6862	)	,
(	6860	)	,
(	6859	)	,
(	6857	)	,
(	6856	)	,
(	6854	)	,
(	6852	)	,
(	6851	)	,
(	6849	)	,
(	6847	)	,
(	6846	)	,
(	6844	)	,
(	6843	)	,
(	6841	)	,
(	6839	)	,
(	6838	)	,
(	6836	)	,
(	6835	)	,
(	6833	)	,
(	6831	)	,
(	6830	)	,
(	6828	)	,
(	6826	)	,
(	6825	)	,
(	6823	)	,
(	6822	)	,
(	6820	)	,
(	6818	)	,
(	6817	)	,
(	6815	)	,
(	6813	)	,
(	6812	)	,
(	6810	)	,
(	6809	)	,
(	6807	)	,
(	6805	)	,
(	6804	)	,
(	6802	)	,
(	6800	)	,
(	6799	)	,
(	6797	)	,
(	6796	)	,
(	6794	)	,
(	6792	)	,
(	6791	)	,
(	6789	)	,
(	6788	)	,
(	6786	)	,
(	6784	)	,
(	6783	)	,
(	6781	)	,
(	6779	)	,
(	6778	)	,
(	6776	)	,
(	6775	)	,
(	6773	)	,
(	6771	)	,
(	6770	)	,
(	6768	)	,
(	6766	)	,
(	6765	)	,
(	6763	)	,
(	6762	)	,
(	6760	)	,
(	6758	)	,
(	6757	)	,
(	6755	)	,
(	6754	)	,
(	6752	)	,
(	6750	)	,
(	6749	)	,
(	6747	)	,
(	6745	)	,
(	6744	)	,
(	6742	)	,
(	6741	)	,
(	6739	)	,
(	6737	)	,
(	6736	)	,
(	6734	)	,
(	6732	)	,
(	6731	)	,
(	6729	)	,
(	6728	)	,
(	6726	)	,
(	6724	)	,
(	6723	)	,
(	6721	)	,
(	6719	)	,
(	6718	)	,
(	6716	)	,
(	6715	)	,
(	6713	)	,
(	6711	)	,
(	6710	)	,
(	6708	)	,
(	6707	)	,
(	6705	)	,
(	6703	)	,
(	6702	)	,
(	6700	)	,
(	6698	)	,
(	6697	)	,
(	6695	)	,
(	6694	)	,
(	6692	)	,
(	6690	)	,
(	6689	)	,
(	6687	)	,
(	6685	)	,
(	6684	)	,
(	6682	)	,
(	6681	)	,
(	6679	)	,
(	6677	)	,
(	6676	)	,
(	6674	)	,
(	6673	)	,
(	6671	)	,
(	6669	)	,
(	6668	)	,
(	6666	)	,
(	6664	)	,
(	6663	)	,
(	6661	)	,
(	6660	)	,
(	6658	)	,
(	6656	)	,
(	6655	)	,
(	6653	)	,
(	6651	)	,
(	6650	)	,
(	6648	)	,
(	6647	)	,
(	6645	)	,
(	6643	)	,
(	6642	)	,
(	6640	)	,
(	6638	)	,
(	6637	)	,
(	6635	)	,
(	6634	)	,
(	6632	)	,
(	6630	)	,
(	6629	)	,
(	6627	)	,
(	6626	)	,
(	6624	)	,
(	6622	)	,
(	6621	)	,
(	6619	)	,
(	6617	)	,
(	6616	)	,
(	6614	)	,
(	6613	)	,
(	6611	)	,
(	6609	)	,
(	6608	)	,
(	6606	)	,
(	6604	)	,
(	6603	)	,
(	6601	)	,
(	6600	)	,
(	6598	)	,
(	6596	)	,
(	6595	)	,
(	6593	)	,
(	6592	)	,
(	6590	)	,
(	6588	)	,
(	6587	)	,
(	6585	)	,
(	6583	)	,
(	6582	)	,
(	6580	)	,
(	6579	)	,
(	6577	)	,
(	6575	)	,
(	6574	)	,
(	6572	)	,
(	6570	)	,
(	6569	)	,
(	6567	)	,
(	6566	)	,
(	6564	)	,
(	6562	)	,
(	6561	)	,
(	6559	)	,
(	6557	)	,
(	6556	)	,
(	6554	)	,
(	6553	)	,
(	6551	)	,
(	6549	)	,
(	6548	)	,
(	6546	)	,
(	6545	)	,
(	6543	)	,
(	6541	)	,
(	6540	)	,
(	6538	)	,
(	6536	)	,
(	6535	)	,
(	6533	)	,
(	6532	)	,
(	6530	)	,
(	6528	)	,
(	6527	)	,
(	6525	)	,
(	6523	)	,
(	6522	)	,
(	6520	)	,
(	6519	)	,
(	6517	)	,
(	6515	)	,
(	6514	)	,
(	6512	)	,
(	6511	)	,
(	6509	)	,
(	6507	)	,
(	6506	)	,
(	6504	)	,
(	6502	)	,
(	6501	)	,
(	6499	)	,
(	6498	)	,
(	6496	)	,
(	6494	)	,
(	6493	)	,
(	6491	)	,
(	6489	)	,
(	6488	)	,
(	6486	)	,
(	6485	)	,
(	6483	)	,
(	6481	)	,
(	6480	)	,
(	6478	)	,
(	6476	)	,
(	6475	)	,
(	6473	)	,
(	6472	)	,
(	6470	)	,
(	6468	)	,
(	6467	)	,
(	6465	)	,
(	6464	)	,
(	6462	)	,
(	6460	)	,
(	6459	)	,
(	6457	)	,
(	6455	)	,
(	6454	)	,
(	6452	)	,
(	6451	)	,
(	6449	)	,
(	6447	)	,
(	6446	)	,
(	6444	)	,
(	6442	)	,
(	6441	)	,
(	6439	)	,
(	6438	)	,
(	6436	)	,
(	6434	)	,
(	6433	)	,
(	6431	)	,
(	6430	)	,
(	6428	)	,
(	6426	)	,
(	6425	)	,
(	6423	)	,
(	6421	)	,
(	6420	)	,
(	6418	)	,
(	6417	)	,
(	6415	)	,
(	6413	)	,
(	6412	)	,
(	6410	)	,
(	6408	)	,
(	6407	)	,
(	6405	)	,
(	6404	)	,
(	6402	)	,
(	6400	)	,
(	6399	)	,
(	6397	)	,
(	6395	)	,
(	6394	)	,
(	6392	)	,
(	6391	)	,
(	6389	)	,
(	6387	)	,
(	6386	)	,
(	6384	)	,
(	6383	)	,
(	6381	)	,
(	6379	)	,
(	6378	)	,
(	6376	)	,
(	6374	)	,
(	6373	)	,
(	6371	)	,
(	6370	)	,
(	6368	)	,
(	6366	)	,
(	6365	)	,
(	6363	)	,
(	6361	)	,
(	6360	)	,
(	6358	)	,
(	6357	)	,
(	6355	)	,
(	6353	)	,
(	6352	)	,
(	6350	)	,
(	6349	)	,
(	6347	)	,
(	6345	)	,
(	6344	)	,
(	6342	)	,
(	6340	)	,
(	6339	)	,
(	6337	)	,
(	6336	)	,
(	6334	)	,
(	6332	)	,
(	6331	)	,
(	6329	)	,
(	6327	)	,
(	6326	)	,
(	6324	)	,
(	6323	)	,
(	6321	)	,
(	6319	)	,
(	6318	)	,
(	6316	)	,
(	6314	)	,
(	6313	)	,
(	6311	)	,
(	6310	)	,
(	6308	)	,
(	6306	)	,
(	6305	)	,
(	6303	)	,
(	6302	)	,
(	6300	)	,
(	6298	)	,
(	6297	)	,
(	6295	)	,
(	6293	)	,
(	6292	)	,
(	6290	)	,
(	6289	)	,
(	6287	)	,
(	6285	)	,
(	6284	)	,
(	6282	)	,
(	6280	)	,
(	6279	)	,
(	6277	)	,
(	6276	)	,
(	6274	)	,
(	6272	)	,
(	6271	)	,
(	6269	)	,
(	6268	)	,
(	6266	)	,
(	6264	)	,
(	6263	)	,
(	6261	)	,
(	6259	)	,
(	6258	)	,
(	6256	)	,
(	6255	)	,
(	6253	)	,
(	6251	)	,
(	6250	)	,
(	6248	)	,
(	6246	)	,
(	6245	)	,
(	6243	)	,
(	6242	)	,
(	6240	)	,
(	6238	)	,
(	6237	)	,
(	6235	)	,
(	6233	)	,
(	6232	)	,
(	6230	)	,
(	6229	)	,
(	6227	)	,
(	6225	)	,
(	6224	)	,
(	6222	)	,
(	6221	)	,
(	6219	)	,
(	6217	)	,
(	6216	)	,
(	6214	)	,
(	6212	)	,
(	6211	)	,
(	6209	)	,
(	6208	)	,
(	6206	)	,
(	6204	)	,
(	6203	)	,
(	6201	)	,
(	6199	)	,
(	6198	)	,
(	6196	)	,
(	6195	)	,
(	6193	)	,
(	6191	)	,
(	6190	)	,
(	6188	)	,
(	6187	)	,
(	6185	)	,
(	6183	)	,
(	6182	)	,
(	6180	)	,
(	6178	)	,
(	6177	)	,
(	6175	)	,
(	6174	)	,
(	6172	)	,
(	6170	)	,
(	6169	)	,
(	6167	)	,
(	6165	)	,
(	6164	)	,
(	6162	)	,
(	6161	)	,
(	6159	)	,
(	6157	)	,
(	6156	)	,
(	6154	)	,
(	6152	)	,
(	6151	)	,
(	6149	)	,
(	6148	)	,
(	6146	)	,
(	6144	)	,
(	6143	)	,
(	6141	)	,
(	6140	)	,
(	6138	)	,
(	6136	)	,
(	6135	)	,
(	6133	)	,
(	6131	)	,
(	6130	)	,
(	6128	)	,
(	6127	)	,
(	6125	)	,
(	6123	)	,
(	6122	)	,
(	6120	)	,
(	6118	)	,
(	6117	)	,
(	6115	)	,
(	6114	)	,
(	6112	)	,
(	6110	)	,
(	6109	)	,
(	6107	)	,
(	6106	)	,
(	6104	)	,
(	6102	)	,
(	6101	)	,
(	6099	)	,
(	6097	)	,
(	6096	)	,
(	6094	)	,
(	6093	)	,
(	6091	)	,
(	6089	)	,
(	6088	)	,
(	6086	)	,
(	6084	)	,
(	6083	)	,
(	6081	)	,
(	6080	)	,
(	6078	)	,
(	6076	)	,
(	6075	)	,
(	6073	)	,
(	6071	)	,
(	6070	)	,
(	6068	)	,
(	6067	)	,
(	6065	)	,
(	6063	)	,
(	6062	)	,
(	6060	)	,
(	6059	)	,
(	6057	)	,
(	6055	)	,
(	6054	)	,
(	6052	)	,
(	6050	)	,
(	6049	)	,
(	6047	)	,
(	6046	)	,
(	6044	)	,
(	6042	)	,
(	6041	)	,
(	6039	)	,
(	6037	)	,
(	6036	)	,
(	6034	)	,
(	6033	)	,
(	6031	)	,
(	6029	)	,
(	6028	)	,
(	6026	)	,
(	6025	)	,
(	6023	)	,
(	6021	)	,
(	6020	)	,
(	6018	)	,
(	6016	)	,
(	6015	)	,
(	6013	)	,
(	6012	)	,
(	6010	)	,
(	6008	)	,
(	6007	)	,
(	6005	)	,
(	6003	)	,
(	6002	)	,
(	6000	)	,
(	5999	)	,
(	5997	)	,
(	5995	)	,
(	5994	)	,
(	5992	)	,
(	5990	)	,
(	5989	)	,
(	5987	)	,
(	5986	)	,
(	5984	)	,
(	5982	)	,
(	5981	)	,
(	5979	)	,
(	5978	)	,
(	5976	)	,
(	5974	)	,
(	5973	)	,
(	5971	)	,
(	5969	)	,
(	5968	)	,
(	5966	)	,
(	5965	)	,
(	5963	)	,
(	5961	)	,
(	5960	)	,
(	5958	)	,
(	5956	)	,
(	5955	)	,
(	5953	)	,
(	5952	)	,
(	5950	)	,
(	5948	)	,
(	5947	)	,
(	5945	)	,
(	5944	)	,
(	5942	)	,
(	5940	)	,
(	5939	)	,
(	5937	)	,
(	5935	)	,
(	5934	)	,
(	5932	)	,
(	5931	)	,
(	5929	)	,
(	5927	)	,
(	5926	)	,
(	5924	)	,
(	5922	)	,
(	5921	)	,
(	5919	)	,
(	5918	)	,
(	5916	)	,
(	5914	)	,
(	5913	)	,
(	5911	)	,
(	5909	)	,
(	5908	)	,
(	5906	)	,
(	5905	)	,
(	5903	)	,
(	5901	)	,
(	5900	)	,
(	5898	)	,
(	5897	)	,
(	5895	)	,
(	5893	)	,
(	5892	)	,
(	5890	)	,
(	5888	)	,
(	5887	)	,
(	5885	)	,
(	5884	)	,
(	5882	)	,
(	5880	)	,
(	5879	)	,
(	5877	)	,
(	5875	)	,
(	5874	)	,
(	5872	)	,
(	5871	)	,
(	5869	)	,
(	5867	)	,
(	5866	)	,
(	5864	)	,
(	5863	)	,
(	5861	)	,
(	5859	)	,
(	5858	)	,
(	5856	)	,
(	5854	)	,
(	5853	)	,
(	5851	)	,
(	5850	)	,
(	5848	)	,
(	5846	)	,
(	5845	)	,
(	5843	)	,
(	5841	)	,
(	5840	)	,
(	5838	)	,
(	5837	)	,
(	5835	)	,
(	5833	)	,
(	5832	)	,
(	5830	)	,
(	5828	)	,
(	5827	)	,
(	5825	)	,
(	5824	)	,
(	5822	)	,
(	5820	)	,
(	5819	)	,
(	5817	)	,
(	5816	)	,
(	5814	)	,
(	5812	)	,
(	5811	)	,
(	5809	)	,
(	5807	)	,
(	5806	)	,
(	5804	)	,
(	5803	)	,
(	5801	)	,
(	5799	)	,
(	5798	)	,
(	5796	)	,
(	5794	)	,
(	5793	)	,
(	5791	)	,
(	5790	)	,
(	5788	)	,
(	5786	)	,
(	5785	)	,
(	5783	)	,
(	5782	)	,
(	5780	)	,
(	5778	)	,
(	5777	)	,
(	5775	)	,
(	5773	)	,
(	5772	)	,
(	5770	)	,
(	5769	)	,
(	5767	)	,
(	5765	)	,
(	5764	)	,
(	5762	)	,
(	5760	)	,
(	5759	)	,
(	5757	)	,
(	5756	)	,
(	5754	)	,
(	5752	)	,
(	5751	)	,
(	5749	)	,
(	5747	)	,
(	5746	)	,
(	5744	)	,
(	5743	)	,
(	5741	)	,
(	5739	)	,
(	5738	)	,
(	5736	)	,
(	5735	)	,
(	5733	)	,
(	5731	)	,
(	5730	)	,
(	5728	)	,
(	5726	)	,
(	5725	)	,
(	5723	)	,
(	5722	)	,
(	5720	)	,
(	5718	)	,
(	5717	)	,
(	5715	)	,
(	5713	)	,
(	5712	)	,
(	5710	)	,
(	5709	)	,
(	5707	)	,
(	5705	)	,
(	5704	)	,
(	5702	)	,
(	5701	)	,
(	5699	)	,
(	5697	)	,
(	5696	)	,
(	5694	)	,
(	5692	)	,
(	5691	)	,
(	5689	)	,
(	5688	)	,
(	5686	)	,
(	5684	)	,
(	5683	)	,
(	5681	)	,
(	5679	)	,
(	5678	)	,
(	5676	)	,
(	5675	)	,
(	5673	)	,
(	5671	)	,
(	5670	)	,
(	5668	)	,
(	5666	)	,
(	5665	)	,
(	5663	)	,
(	5662	)	,
(	5660	)	,
(	5658	)	,
(	5657	)	,
(	5655	)	,
(	5654	)	,
(	5652	)	,
(	5650	)	,
(	5649	)	,
(	5647	)	,
(	5645	)	,
(	5644	)	,
(	5642	)	,
(	5641	)	,
(	5639	)	,
(	5637	)	,
(	5636	)	,
(	5634	)	,
(	5632	)	,
(	5631	)	,
(	5629	)	,
(	5628	)	,
(	5626	)	,
(	5624	)	,
(	5623	)	,
(	5621	)	,
(	5620	)	,
(	5618	)	,
(	5616	)	,
(	5615	)	,
(	5613	)	,
(	5611	)	,
(	5610	)	,
(	5608	)	,
(	5607	)	,
(	5605	)	,
(	5603	)	,
(	5602	)	,
(	5600	)	,
(	5598	)	,
(	5597	)	,
(	5595	)	,
(	5594	)	,
(	5592	)	,
(	5590	)	,
(	5589	)	,
(	5587	)	,
(	5585	)	,
(	5584	)	,
(	5582	)	,
(	5581	)	,
(	5579	)	,
(	5577	)	,
(	5576	)	,
(	5574	)	,
(	5573	)	,
(	5571	)	,
(	5569	)	,
(	5568	)	,
(	5566	)	,
(	5564	)	,
(	5563	)	,
(	5561	)	,
(	5560	)	,
(	5558	)	,
(	5556	)	,
(	5555	)	,
(	5553	)	,
(	5551	)	,
(	5550	)	,
(	5548	)	,
(	5547	)	,
(	5545	)	,
(	5543	)	,
(	5542	)	,
(	5540	)	,
(	5539	)	,
(	5537	)	,
(	5535	)	,
(	5534	)	,
(	5532	)	,
(	5530	)	,
(	5529	)	,
(	5527	)	,
(	5526	)	,
(	5524	)	,
(	5522	)	,
(	5521	)	,
(	5519	)	,
(	5517	)	,
(	5516	)	,
(	5514	)	,
(	5513	)	,
(	5511	)	,
(	5509	)	,
(	5508	)	,
(	5506	)	,
(	5504	)	,
(	5503	)	,
(	5501	)	,
(	5500	)	,
(	5498	)	,
(	5496	)	,
(	5495	)	,
(	5493	)	,
(	5492	)	,
(	5490	)	,
(	5488	)	,
(	5487	)	,
(	5485	)	,
(	5483	)	,
(	5482	)	,
(	5480	)	,
(	5479	)	,
(	5477	)	,
(	5475	)	,
(	5474	)	,
(	5472	)	,
(	5470	)	,
(	5469	)	,
(	5467	)	,
(	5466	)	,
(	5464	)	,
(	5462	)	,
(	5461	)	,
(	5459	)	,
(	5458	)	,
(	5456	)	,
(	5454	)	,
(	5453	)	,
(	5451	)	,
(	5449	)	,
(	5448	)	,
(	5446	)	,
(	5445	)	,
(	5443	)	,
(	5441	)	,
(	5440	)	,
(	5438	)	,
(	5436	)	,
(	5435	)	,
(	5433	)	,
(	5432	)	,
(	5430	)	,
(	5428	)	,
(	5427	)	,
(	5425	)	,
(	5423	)	,
(	5422	)	,
(	5420	)	,
(	5419	)	,
(	5417	)	,
(	5415	)	,
(	5414	)	,
(	5412	)	,
(	5411	)	,
(	5409	)	,
(	5407	)	,
(	5406	)	,
(	5404	)	,
(	5402	)	,
(	5401	)	,
(	5399	)	,
(	5398	)	,
(	5396	)	,
(	5394	)	,
(	5393	)	,
(	5391	)	,
(	5389	)	,
(	5388	)	,
(	5386	)	,
(	5385	)	,
(	5383	)	,
(	5381	)	,
(	5380	)	,
(	5378	)	,
(	5377	)	,
(	5375	)	,
(	5373	)	,
(	5372	)	,
(	5370	)	,
(	5368	)	,
(	5367	)	,
(	5365	)	,
(	5364	)	,
(	5362	)	,
(	5360	)	,
(	5359	)	,
(	5357	)	,
(	5355	)	,
(	5354	)	,
(	5352	)	,
(	5351	)	,
(	5349	)	,
(	5347	)	,
(	5346	)	,
(	5344	)	,
(	5342	)	,
(	5341	)	,
(	5339	)	,
(	5338	)	,
(	5336	)	,
(	5334	)	,
(	5333	)	,
(	5331	)	,
(	5330	)	,
(	5328	)	,
(	5326	)	,
(	5325	)	,
(	5323	)	,
(	5321	)	,
(	5320	)	,
(	5318	)	,
(	5317	)	,
(	5315	)	,
(	5313	)	,
(	5312	)	,
(	5310	)	,
(	5308	)	,
(	5307	)	,
(	5305	)	,
(	5304	)	,
(	5302	)	,
(	5300	)	,
(	5299	)	,
(	5297	)	,
(	5296	)	,
(	5294	)	,
(	5292	)	,
(	5291	)	,
(	5289	)	,
(	5287	)	,
(	5286	)	,
(	5284	)	,
(	5283	)	,
(	5281	)	,
(	5279	)	,
(	5278	)	,
(	5276	)	,
(	5274	)	,
(	5273	)	,
(	5271	)	,
(	5270	)	,
(	5268	)	,
(	5266	)	,
(	5265	)	,
(	5263	)	,
(	5261	)	,
(	5260	)	,
(	5258	)	,
(	5257	)	,
(	5255	)	,
(	5253	)	,
(	5252	)	,
(	5250	)	,
(	5249	)	,
(	5247	)	,
(	5245	)	,
(	5244	)	,
(	5242	)	,
(	5240	)	,
(	5239	)	,
(	5237	)	,
(	5236	)	,
(	5234	)	,
(	5232	)	,
(	5231	)	,
(	5229	)	,
(	5227	)	,
(	5226	)	,
(	5224	)	,
(	5223	)	,
(	5221	)	,
(	5219	)	,
(	5218	)	,
(	5216	)	,
(	5215	)	,
(	5213	)	,
(	5211	)	,
(	5210	)	,
(	5208	)	,
(	5206	)	,
(	5205	)	,
(	5203	)	,
(	5202	)	,
(	5200	)	,
(	5198	)	,
(	5197	)	,
(	5195	)	,
(	5193	)	,
(	5192	)	,
(	5190	)	,
(	5189	)	,
(	5187	)	,
(	5185	)	,
(	5184	)	,
(	5182	)	,
(	5180	)	,
(	5179	)	,
(	5177	)	,
(	5176	)	,
(	5174	)	,
(	5172	)	,
(	5171	)	,
(	5169	)	,
(	5168	)	,
(	5166	)	,
(	5164	)	,
(	5163	)	,
(	5161	)	,
(	5159	)	,
(	5158	)	,
(	5156	)	,
(	5155	)	,
(	5153	)	,
(	5151	)	,
(	5150	)	,
(	5148	)	,
(	5146	)	,
(	5145	)	,
(	5143	)	,
(	5142	)	,
(	5140	)	,
(	5138	)	,
(	5137	)	,
(	5135	)	,
(	5134	)	,
(	5132	)	,
(	5130	)	,
(	5129	)	,
(	5127	)	,
(	5125	)	,
(	5124	)	,
(	5122	)	,
(	5121	)	,
(	5119	)	,
(	5117	)	,
(	5116	)	,
(	5114	)	,
(	5112	)	,
(	5111	)	,
(	5109	)	,
(	5108	)	,
(	5106	)	,
(	5104	)	,
(	5103	)	,
(	5101	)	,
(	5099	)	,
(	5098	)	,
(	5096	)	,
(	5095	)	,
(	5093	)	,
(	5091	)	,
(	5090	)	,
(	5088	)	,
(	5087	)	,
(	5085	)	,
(	5083	)	,
(	5082	)	,
(	5080	)	,
(	5078	)	,
(	5077	)	,
(	5075	)	,
(	5074	)	,
(	5072	)	,
(	5070	)	,
(	5069	)	,
(	5067	)	,
(	5065	)	,
(	5064	)	,
(	5062	)	,
(	5061	)	,
(	5059	)	,
(	5057	)	,
(	5056	)	,
(	5054	)	,
(	5053	)	,
(	5051	)	,
(	5049	)	,
(	5048	)	,
(	5046	)	,
(	5044	)	,
(	5043	)	,
(	5041	)	,
(	5040	)	,
(	5038	)	,
(	5036	)	,
(	5035	)	,
(	5033	)	,
(	5031	)	,
(	5030	)	,
(	5028	)	,
(	5027	)	,
(	5025	)	,
(	5023	)	,
(	5022	)	,
(	5020	)	,
(	5018	)	,
(	5017	)	,
(	5015	)	,
(	5014	)	,
(	5012	)	,
(	5010	)	,
(	5009	)	,
(	5007	)	,
(	5006	)	,
(	5004	)	,
(	5002	)	,
(	5001	)	,
(	4999	)	,
(	4997	)	,
(	4996	)	,
(	4994	)	,
(	4993	)	,
(	4991	)	,
(	4989	)	,
(	4988	)	,
(	4986	)	,
(	4984	)	,
(	4983	)	,
(	4981	)	,
(	4980	)	,
(	4978	)	,
(	4976	)	,
(	4975	)	,
(	4973	)	,
(	4972	)	,
(	4970	)	,
(	4968	)	,
(	4967	)	,
(	4965	)	,
(	4963	)	,
(	4962	)	,
(	4960	)	,
(	4959	)	,
(	4957	)	,
(	4955	)	,
(	4954	)	,
(	4952	)	,
(	4950	)	,
(	4949	)	,
(	4947	)	,
(	4946	)	,
(	4944	)	,
(	4942	)	,
(	4941	)	,
(	4939	)	,
(	4937	)	,
(	4936	)	,
(	4934	)	,
(	4933	)	,
(	4931	)	,
(	4929	)	,
(	4928	)	,
(	4926	)	,
(	4925	)	,
(	4923	)	,
(	4921	)	,
(	4920	)	,
(	4918	)	,
(	4916	)	,
(	4915	)	,
(	4913	)	,
(	4912	)	,
(	4910	)	,
(	4908	)	,
(	4907	)	,
(	4905	)	,
(	4903	)	,
(	4902	)	,
(	4900	)	,
(	4899	)	,
(	4897	)	,
(	4895	)	,
(	4894	)	,
(	4892	)	,
(	4891	)	,
(	4889	)	,
(	4887	)	,
(	4886	)	,
(	4884	)	,
(	4882	)	,
(	4881	)	,
(	4879	)	,
(	4878	)	,
(	4876	)	,
(	4874	)	,
(	4873	)	,
(	4871	)	,
(	4869	)	,
(	4868	)	,
(	4866	)	,
(	4865	)	,
(	4863	)	,
(	4861	)	,
(	4860	)	,
(	4858	)	,
(	4856	)	,
(	4855	)	,
(	4853	)	,
(	4852	)	,
(	4850	)	,
(	4848	)	,
(	4847	)	,
(	4845	)	,
(	4844	)	,
(	4842	)	,
(	4840	)	,
(	4839	)	,
(	4837	)	,
(	4835	)	,
(	4834	)	,
(	4832	)	,
(	4831	)	,
(	4829	)	,
(	4827	)	,
(	4826	)	,
(	4824	)	,
(	4822	)	,
(	4821	)	,
(	4819	)	,
(	4818	)	,
(	4816	)	,
(	4814	)	,
(	4813	)	,
(	4811	)	,
(	4810	)	,
(	4808	)	,
(	4806	)	,
(	4805	)	,
(	4803	)	,
(	4801	)	,
(	4800	)	,
(	4798	)	,
(	4797	)	,
(	4795	)	,
(	4793	)	,
(	4792	)	,
(	4790	)	,
(	4788	)	,
(	4787	)	,
(	4785	)	,
(	4784	)	,
(	4782	)	,
(	4780	)	,
(	4779	)	,
(	4777	)	,
(	4775	)	,
(	4774	)	,
(	4772	)	,
(	4771	)	,
(	4769	)	,
(	4767	)	,
(	4766	)	,
(	4764	)	,
(	4763	)	,
(	4761	)	,
(	4759	)	,
(	4758	)	,
(	4756	)	,
(	4754	)	,
(	4753	)	,
(	4751	)	,
(	4750	)	,
(	4748	)	,
(	4746	)	,
(	4745	)	,
(	4743	)	,
(	4741	)	,
(	4740	)	,
(	4738	)	,
(	4737	)	,
(	4735	)	,
(	4733	)	,
(	4732	)	,
(	4730	)	,
(	4729	)	,
(	4727	)	,
(	4725	)	,
(	4724	)	,
(	4722	)	,
(	4720	)	,
(	4719	)	,
(	4717	)	,
(	4716	)	,
(	4714	)	,
(	4712	)	,
(	4711	)	,
(	4709	)	,
(	4707	)	,
(	4706	)	,
(	4704	)	,
(	4703	)	,
(	4701	)	,
(	4699	)	,
(	4698	)	,
(	4696	)	,
(	4694	)	,
(	4693	)	,
(	4691	)	,
(	4690	)	,
(	4688	)	,
(	4686	)	,
(	4685	)	,
(	4683	)	,
(	4682	)	,
(	4680	)	,
(	4678	)	,
(	4677	)	,
(	4675	)	,
(	4673	)	,
(	4672	)	,
(	4670	)	,
(	4669	)	,
(	4667	)	,
(	4665	)	,
(	4664	)	,
(	4662	)	,
(	4660	)	,
(	4659	)	,
(	4657	)	,
(	4656	)	,
(	4654	)	,
(	4652	)	,
(	4651	)	,
(	4649	)	,
(	4648	)	,
(	4646	)	,
(	4644	)	,
(	4643	)	,
(	4641	)	,
(	4639	)	,
(	4638	)	,
(	4636	)	,
(	4635	)	,
(	4633	)	,
(	4631	)	,
(	4630	)	,
(	4628	)	,
(	4626	)	,
(	4625	)	,
(	4623	)	,
(	4622	)	,
(	4620	)	,
(	4618	)	,
(	4617	)	,
(	4615	)	,
(	4613	)	,
(	4612	)	,
(	4610	)	,
(	4609	)	,
(	4607	)	,
(	4605	)	,
(	4604	)	,
(	4602	)	,
(	4601	)	,
(	4599	)	,
(	4597	)	,
(	4596	)	,
(	4594	)	,
(	4592	)	,
(	4591	)	,
(	4589	)	,
(	4588	)	,
(	4586	)	,
(	4584	)	,
(	4583	)	,
(	4581	)	,
(	4579	)	,
(	4578	)	,
(	4576	)	,
(	4575	)	,
(	4573	)	,
(	4571	)	,
(	4570	)	,
(	4568	)	,
(	4567	)	,
(	4565	)	,
(	4563	)	,
(	4562	)	,
(	4560	)	,
(	4558	)	,
(	4557	)	,
(	4555	)	,
(	4554	)	,
(	4552	)	,
(	4550	)	,
(	4549	)	,
(	4547	)	,
(	4545	)	,
(	4544	)	,
(	4542	)	,
(	4541	)	,
(	4539	)	,
(	4537	)	,
(	4536	)	,
(	4534	)	,
(	4532	)	,
(	4531	)	,
(	4529	)	,
(	4528	)	,
(	4526	)	,
(	4524	)	,
(	4523	)	,
(	4521	)	,
(	4520	)	,
(	4518	)	,
(	4516	)	,
(	4515	)	,
(	4513	)	,
(	4511	)	,
(	4510	)	,
(	4508	)	,
(	4507	)	,
(	4505	)	,
(	4503	)	,
(	4502	)	,
(	4500	)	,
(	4498	)	,
(	4497	)	,
(	4495	)	,
(	4494	)	,
(	4492	)	,
(	4490	)	,
(	4489	)	,
(	4487	)	,
(	4486	)	,
(	4484	)	,
(	4482	)	,
(	4481	)	,
(	4479	)	,
(	4477	)	,
(	4476	)	,
(	4474	)	,
(	4473	)	,
(	4471	)	,
(	4469	)	,
(	4468	)	,
(	4466	)	,
(	4464	)	,
(	4463	)	,
(	4461	)	,
(	4460	)	,
(	4458	)	,
(	4456	)	,
(	4455	)	,
(	4453	)	,
(	4451	)	,
(	4450	)	,
(	4448	)	,
(	4447	)	,
(	4445	)	,
(	4443	)	,
(	4442	)	,
(	4440	)	,
(	4439	)	,
(	4437	)	,
(	4435	)	,
(	4434	)	,
(	4432	)	,
(	4430	)	,
(	4429	)	,
(	4427	)	,
(	4426	)	,
(	4424	)	,
(	4422	)	,
(	4421	)	,
(	4419	)	,
(	4417	)	,
(	4416	)	,
(	4414	)	,
(	4413	)	,
(	4411	)	,
(	4409	)	,
(	4408	)	,
(	4406	)	,
(	4405	)	,
(	4403	)	,
(	4401	)	,
(	4400	)	,
(	4398	)	,
(	4396	)	,
(	4395	)	,
(	4393	)	,
(	4392	)	,
(	4390	)	,
(	4388	)	,
(	4387	)	,
(	4385	)	,
(	4383	)	,
(	4382	)	,
(	4380	)	,
(	4379	)	,
(	4377	)	,
(	4375	)	,
(	4374	)	,
(	4372	)	,
(	4370	)	,
(	4369	)	,
(	4367	)	,
(	4366	)	,
(	4364	)	,
(	4362	)	,
(	4361	)	,
(	4359	)	,
(	4358	)	,
(	4356	)	,
(	4354	)	,
(	4353	)	,
(	4351	)	,
(	4349	)	,
(	4348	)	,
(	4346	)	,
(	4345	)	,
(	4343	)	,
(	4341	)	,
(	4340	)	,
(	4338	)	,
(	4336	)	,
(	4335	)	,
(	4333	)	,
(	4332	)	,
(	4330	)	,
(	4328	)	,
(	4327	)	,
(	4325	)	,
(	4324	)	,
(	4322	)	,
(	4320	)	,
(	4319	)	,
(	4317	)	,
(	4315	)	,
(	4314	)	,
(	4312	)	,
(	4311	)	,
(	4309	)	,
(	4307	)	,
(	4306	)	,
(	4304	)	,
(	4302	)	,
(	4301	)	,
(	4299	)	,
(	4298	)	,
(	4296	)	,
(	4294	)	,
(	4293	)	,
(	4291	)	,
(	4289	)	,
(	4288	)	,
(	4286	)	,
(	4285	)	,
(	4283	)	,
(	4281	)	,
(	4280	)	,
(	4278	)	,
(	4277	)	,
(	4275	)	,
(	4273	)	,
(	4272	)	,
(	4270	)	,
(	4268	)	,
(	4267	)	,
(	4265	)	,
(	4264	)	,
(	4262	)	,
(	4260	)	,
(	4259	)	,
(	4257	)	,
(	4255	)	,
(	4254	)	,
(	4252	)	,
(	4251	)	,
(	4249	)	,
(	4247	)	,
(	4246	)	,
(	4244	)	,
(	4243	)	,
(	4241	)	,
(	4239	)	,
(	4238	)	,
(	4236	)	,
(	4234	)	,
(	4233	)	,
(	4231	)	,
(	4230	)	,
(	4228	)	,
(	4226	)	,
(	4225	)	,
(	4223	)	,
(	4221	)	,
(	4220	)	,
(	4218	)	,
(	4217	)	,
(	4215	)	,
(	4213	)	,
(	4212	)	,
(	4210	)	,
(	4208	)	,
(	4207	)	,
(	4205	)	,
(	4204	)	,
(	4202	)	,
(	4200	)	,
(	4199	)	,
(	4197	)	,
(	4196	)	,
(	4194	)	,
(	4192	)	,
(	4191	)	,
(	4189	)	,
(	4187	)	,
(	4186	)	,
(	4184	)	,
(	4183	)	,
(	4181	)	,
(	4179	)	,
(	4178	)	,
(	4176	)	,
(	4174	)	,
(	4173	)	,
(	4171	)	,
(	4170	)	,
(	4168	)	,
(	4166	)	,
(	4165	)	,
(	4163	)	,
(	4162	)	,
(	4160	)	,
(	4158	)	,
(	4157	)	,
(	4155	)	,
(	4153	)	,
(	4152	)	,
(	4150	)	,
(	4149	)	,
(	4147	)	,
(	4145	)	,
(	4144	)	,
(	4142	)	,
(	4140	)	,
(	4139	)	,
(	4137	)	,
(	4136	)	,
(	4134	)	,
(	4132	)	,
(	4131	)	,
(	4129	)	,
(	4127	)	,
(	4126	)	,
(	4124	)	,
(	4123	)	,
(	4121	)	,
(	4119	)	,
(	4118	)	,
(	4116	)	,
(	4115	)	,
(	4113	)	,
(	4111	)	,
(	4110	)	,
(	4108	)	,
(	4106	)	,
(	4105	)	,
(	4103	)	,
(	4102	)	,
(	4100	)	,
(	4098	)	,
(	4097	)	,
(	4095	)	,
(	4093	)	,
(	4092	)	,
(	4090	)	,
(	4089	)	,
(	4087	)	,
(	4085	)	,
(	4084	)	,
(	4082	)	,
(	4081	)	,
(	4079	)	,
(	4077	)	,
(	4076	)	,
(	4074	)	,
(	4072	)	,
(	4071	)	,
(	4069	)	,
(	4068	)	,
(	4066	)	,
(	4064	)	,
(	4063	)	,
(	4061	)	,
(	4059	)	,
(	4058	)	,
(	4056	)	,
(	4055	)	,
(	4053	)	,
(	4051	)	,
(	4050	)	,
(	4048	)	,
(	4046	)	,
(	4045	)	,
(	4043	)	,
(	4042	)	,
(	4040	)	,
(	4038	)	,
(	4037	)	,
(	4035	)	,
(	4034	)	,
(	4032	)	,
(	4030	)	,
(	4029	)	,
(	4027	)	,
(	4025	)	,
(	4024	)	,
(	4022	)	,
(	4021	)	,
(	4019	)	,
(	4017	)	,
(	4016	)	,
(	4014	)	,
(	4012	)	,
(	4011	)	,
(	4009	)	,
(	4008	)	,
(	4006	)	,
(	4004	)	,
(	4003	)	,
(	4001	)	,
(	4000	)	,
(	3998	)	,
(	3996	)	,
(	3995	)	,
(	3993	)	,
(	3991	)	,
(	3990	)	,
(	3988	)	,
(	3987	)	,
(	3985	)	,
(	3983	)	,
(	3982	)	,
(	3980	)	,
(	3978	)	,
(	3977	)	,
(	3975	)	,
(	3974	)	,
(	3972	)	,
(	3970	)	,
(	3969	)	,
(	3967	)	,
(	3965	)	,
(	3964	)	,
(	3962	)	,
(	3961	)	,
(	3959	)	,
(	3957	)	,
(	3956	)	,
(	3954	)	,
(	3953	)	,
(	3951	)	,
(	3949	)	,
(	3948	)	,
(	3946	)	,
(	3944	)	,
(	3943	)	,
(	3941	)	,
(	3940	)	,
(	3938	)	,
(	3936	)	,
(	3935	)	,
(	3933	)	,
(	3931	)	,
(	3930	)	,
(	3928	)	,
(	3927	)	,
(	3925	)	,
(	3923	)	,
(	3922	)	,
(	3920	)	,
(	3919	)	,
(	3917	)	,
(	3915	)	,
(	3914	)	,
(	3912	)	,
(	3910	)	,
(	3909	)	,
(	3907	)	,
(	3906	)	,
(	3904	)	,
(	3902	)	,
(	3901	)	,
(	3899	)	,
(	3897	)	,
(	3896	)	,
(	3894	)	,
(	3893	)	,
(	3891	)	,
(	3889	)	,
(	3888	)	,
(	3886	)	,
(	3884	)	,
(	3883	)	,
(	3881	)	,
(	3880	)	,
(	3878	)	,
(	3876	)	,
(	3875	)	,
(	3873	)	,
(	3872	)	,
(	3870	)	,
(	3868	)	,
(	3867	)	,
(	3865	)	,
(	3863	)	,
(	3862	)	,
(	3860	)	,
(	3859	)	,
(	3857	)	,
(	3855	)	,
(	3854	)	,
(	3852	)	,
(	3850	)	,
(	3849	)	,
(	3847	)	,
(	3846	)	,
(	3844	)	,
(	3842	)	,
(	3841	)	,
(	3839	)	,
(	3838	)	,
(	3836	)	,
(	3834	)	,
(	3833	)	,
(	3831	)	,
(	3829	)	,
(	3828	)	,
(	3826	)	,
(	3825	)	,
(	3823	)	,
(	3821	)	,
(	3820	)	,
(	3818	)	,
(	3816	)	,
(	3815	)	,
(	3813	)	,
(	3812	)	,
(	3810	)	,
(	3808	)	,
(	3807	)	,
(	3805	)	,
(	3803	)	,
(	3802	)	,
(	3800	)	,
(	3799	)	,
(	3797	)	,
(	3795	)	,
(	3794	)	,
(	3792	)	,
(	3791	)	,
(	3789	)	,
(	3787	)	,
(	3786	)	,
(	3784	)	,
(	3782	)	,
(	3781	)	,
(	3779	)	,
(	3778	)	,
(	3776	)	,
(	3774	)	,
(	3773	)	,
(	3771	)	,
(	3769	)	,
(	3768	)	,
(	3766	)	,
(	3765	)	,
(	3763	)	,
(	3761	)	,
(	3760	)	,
(	3758	)	,
(	3757	)	,
(	3755	)	,
(	3753	)	,
(	3752	)	,
(	3750	)	,
(	3748	)	,
(	3747	)	,
(	3745	)	,
(	3744	)	,
(	3742	)	,
(	3740	)	,
(	3739	)	,
(	3737	)	,
(	3735	)	,
(	3734	)	,
(	3732	)	,
(	3731	)	,
(	3729	)	,
(	3727	)	,
(	3726	)	,
(	3724	)	,
(	3722	)	,
(	3721	)	,
(	3719	)	,
(	3718	)	,
(	3716	)	,
(	3714	)	,
(	3713	)	,
(	3711	)	,
(	3710	)	,
(	3708	)	,
(	3706	)	,
(	3705	)	,
(	3703	)	,
(	3701	)	,
(	3700	)	,
(	3698	)	,
(	3697	)	,
(	3695	)	,
(	3693	)	,
(	3692	)	,
(	3690	)	,
(	3688	)	,
(	3687	)	,
(	3685	)	,
(	3684	)	,
(	3682	)	,
(	3680	)	,
(	3679	)	,
(	3677	)	,
(	3676	)	,
(	3674	)	,
(	3672	)	,
(	3671	)	,
(	3669	)	,
(	3667	)	,
(	3666	)	,
(	3664	)	,
(	3663	)	,
(	3661	)	,
(	3659	)	,
(	3658	)	,
(	3656	)	,
(	3654	)	,
(	3653	)	,
(	3651	)	,
(	3650	)	,
(	3648	)	,
(	3646	)	,
(	3645	)	,
(	3643	)	,
(	3641	)	,
(	3640	)	,
(	3638	)	,
(	3637	)	,
(	3635	)	,
(	3633	)	,
(	3632	)	,
(	3630	)	,
(	3629	)	,
(	3627	)	,
(	3625	)	,
(	3624	)	,
(	3622	)	,
(	3620	)	,
(	3619	)	,
(	3617	)	,
(	3616	)	,
(	3614	)	,
(	3612	)	,
(	3611	)	,
(	3609	)	,
(	3607	)	,
(	3606	)	,
(	3604	)	,
(	3603	)	,
(	3601	)	,
(	3599	)	,
(	3598	)	,
(	3596	)	,
(	3595	)	,
(	3593	)	,
(	3591	)	,
(	3590	)	,
(	3588	)	,
(	3586	)	,
(	3585	)	,
(	3583	)	,
(	3582	)	,
(	3580	)	,
(	3578	)	,
(	3577	)	,
(	3575	)	,
(	3573	)	,
(	3572	)	,
(	3570	)	,
(	3569	)	,
(	3567	)	,
(	3565	)	,
(	3564	)	,
(	3562	)	,
(	3560	)	,
(	3559	)	,
(	3557	)	,
(	3556	)	,
(	3554	)	,
(	3552	)	,
(	3551	)	,
(	3549	)	,
(	3548	)	,
(	3546	)	,
(	3544	)	,
(	3543	)	,
(	3541	)	,
(	3539	)	,
(	3538	)	,
(	3536	)	,
(	3535	)	,
(	3533	)	,
(	3531	)	,
(	3530	)	,
(	3528	)	,
(	3526	)	,
(	3525	)	,
(	3523	)	,
(	3522	)	,
(	3520	)	,
(	3518	)	,
(	3517	)	,
(	3515	)	,
(	3514	)	,
(	3512	)	,
(	3510	)	,
(	3509	)	,
(	3507	)	,
(	3505	)	,
(	3504	)	,
(	3502	)	,
(	3501	)	,
(	3499	)	,
(	3497	)	,
(	3496	)	,
(	3494	)	,
(	3492	)	,
(	3491	)	,
(	3489	)	,
(	3488	)	,
(	3486	)	,
(	3484	)	,
(	3483	)	,
(	3481	)	,
(	3479	)	,
(	3478	)	,
(	3476	)	,
(	3475	)	,
(	3473	)	,
(	3471	)	,
(	3470	)	,
(	3468	)	,
(	3467	)	,
(	3465	)	,
(	3463	)	,
(	3462	)	,
(	3460	)	,
(	3458	)	,
(	3457	)	,
(	3455	)	,
(	3454	)	,
(	3452	)	,
(	3450	)	,
(	3449	)	,
(	3447	)	,
(	3445	)	,
(	3444	)	,
(	3442	)	,
(	3441	)	,
(	3439	)	,
(	3437	)	,
(	3436	)	,
(	3434	)	,
(	3433	)	,
(	3431	)	,
(	3429	)	,
(	3428	)	,
(	3426	)	,
(	3424	)	,
(	3423	)	,
(	3421	)	,
(	3420	)	,
(	3418	)	,
(	3416	)	,
(	3415	)	,
(	3413	)	,
(	3411	)	,
(	3410	)	,
(	3408	)	,
(	3407	)	,
(	3405	)	,
(	3403	)	,
(	3402	)	,
(	3400	)	,
(	3398	)	,
(	3397	)	,
(	3395	)	,
(	3394	)	,
(	3392	)	,
(	3390	)	,
(	3389	)	,
(	3387	)	,
(	3386	)	,
(	3384	)	,
(	3382	)	,
(	3381	)	,
(	3379	)	,
(	3377	)	,
(	3376	)	,
(	3374	)	,
(	3373	)	,
(	3371	)	,
(	3369	)	,
(	3368	)	,
(	3366	)		-- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the distance input in the v2f_LUT look-up table, and outputs the 
	-- frequency (max counter value for the PWM).
    	
   frequency <= v2f_LUT(to_integer(unsigned(voltage)));

end behavior;
